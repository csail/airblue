../../parameters/WiFi/Macros.bsv