/////////////////////////////////////////////////////////////////////////
// Macros definitions
////////////////////////////////////////////////////////////////////////

// if this SoftPhyHints is defined, we are going to expose it to the external interface
//`define SOFT_PHY_HINTS 1