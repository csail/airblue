//*************************************************************
// Type definitions for use in the Reed-Solomon modules
//-------------------------------------------------------------


// Byte	primitive_polynomial = 8'b00011101;
typedef Bit#(8)   Polynomial;
typedef Bit#(8)	Byte;
typedef Bit#(16)  Word;
