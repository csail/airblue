// total ber: 0.006535
// a = 0.640000 b = 0.000000
// generated by compute-ber.py
// table for rate 0 (curve fit)
// (computed without odd hints)

import Real::*;

function data_t get_ber_r0_log(Bit#(8) hint)
      provisos (RealLiteral#(data_t), Arith#(data_t));
   case (hint) matches
       0: return -1.000000000000000;
       1: return -1.534301141300769;
       2: return -2.200579595346998;
       3: return -2.967345422642400;
       4: return -3.800725711789279;
       5: return -4.674264606465106;
       6: return -5.570629124044506;
       7: return -6.479532481913688;
       8: return -7.395194528746716;
       9: return -8.314462380984828;
      10: return -9.235643392854302;
      11: return -10.157836517923325;
      12: return -11.080564249019554;
      13: return -12.003574131944424;
      14: return -12.926732863238305;
      15: return -13.849970101137506;
      16: return -14.773248740534070;
      17: return -15.696549212172435;
      18: return -16.619861196216359;
      19: return -17.543179250784039;
      20: return -18.466500506326131;
      21: return -19.389823449727029;
      22: return -20.313147283125652;
      23: return -21.236471585814051;
      24: return -22.159796135955585;
      25: return -23.083120816577345;
      26: return -24.006445566000355;
      27: return -24.929770351701741;
      28: return -25.853095156532444;
      29: return -26.776419971449887;
      30: return -27.699744791686001;
      31: return -28.623069614726607;
      32: return -29.546394439245994;
      33: return -30.469719264545144;
      34: return -31.393044090255440;
      35: return -32.316368916182540;
      36: return -33.239693742223956;
      37: return -34.163018568325654;
      38: return -35.086343394459142;
      39: return -36.009668220609385;
      40: return -36.932993046768459;
      41: return -37.856317872932202;
      42: return -38.779642699098389;
      43: return -39.702967525265883;
      44: return -40.626292351434060;
      45: return -41.549617177602592;
      46: return -42.472942003771323;
      47: return -43.396266829940146;
      48: return -44.319591656109026;
      49: return -45.242916482277927;
      50: return -46.166241308446850;
      51: return -47.089566134615779;
      52: return -48.012890960784702;
      53: return -48.936215786953646;
      54: return -49.859540613122583;
      55: return -50.782865439291520;
      56: return -51.706190265460457;
      57: return -52.629515091629393;
      58: return -53.552839917798323;
      59: return -54.476164743967260;
      60: return -55.399489570136197;
      61: return -56.322814396305134;
      62: return -57.246139222474071;
      63: return -58.169464048643007;
      default: return -63;
   endcase
endfunction
