// generated by compute-ber.py
// table for rate 5 (exact)
// (computed without odd hints)

import Real::*;

function data_t get_ber_r5_log(Bit#(8) hint)
      provisos (RealLiteral#(data_t), Arith#(data_t));
   case (hint) matches
       0: return -1.000000000000000;
       1: return -1.357982966361119;
       2: return -1.832908043822234;
       3: return -2.268302648524245;
       4: return -2.959769950744311;
       5: return -3.391337446776092;
       6: return -4.289097956471079;
       7: return -4.615147756280005;
       8: return -5.781889073695585;
       9: return -5.883537520130624;
      10: return -7.373502260908706;
      11: return -7.213941518985686;
      12: return -9.047397162699419;
      13: return -8.543784061780668;
      14: return -10.762907319503853;
      15: return -9.822768710542936;
      16: return -12.505372946201600;
      17: return -11.072512807945250;
      18: return -14.295055381728492;
      19: return -12.242056426678587;
      20: return -15.990225369967208;
      21: return -14.066972402299101;
      22: return -17.734433351337639;
      23: return -14.737241473820978;
      24: return -19.398274718961950;
      25: return -18.029324976419364;
      26: return -21.706790226648341;
      27: return -63.000000000000000;
      28: return -23.596159683605332;
      29: return -63.000000000000000;
      30: return -63.000000000000000;
      31: return -63.000000000000000;
      32: return -63.000000000000000;
      33: return -63.000000000000000;
      34: return -63.000000000000000;
      35: return -63.000000000000000;
      36: return -63.000000000000000;
      37: return -63.000000000000000;
      38: return -63.000000000000000;
      39: return -63.000000000000000;
      40: return -63.000000000000000;
      41: return -63.000000000000000;
      42: return -63.000000000000000;
      43: return -63.000000000000000;
      44: return -63.000000000000000;
      45: return -63.000000000000000;
      46: return -63.000000000000000;
      47: return -63.000000000000000;
      48: return -63.000000000000000;
      49: return -63.000000000000000;
      50: return -63.000000000000000;
      51: return -63.000000000000000;
      52: return -63.000000000000000;
      53: return -63.000000000000000;
      54: return -63.000000000000000;
      55: return -63.000000000000000;
      56: return -63.000000000000000;
      57: return -63.000000000000000;
      58: return -63.000000000000000;
      59: return -63.000000000000000;
      60: return -63.000000000000000;
      61: return -63.000000000000000;
      62: return -63.000000000000000;
      63: return -63.000000000000000;
      default: return -63;
   endcase
endfunction
