// generated by compute-ber.py
// table for rate 1 (exact)
// (computed without odd hints)

import Real::*;

function data_t get_ber_r1_log(Bit#(8) hint)
      provisos (RealLiteral#(data_t), Arith#(data_t));
   case (hint) matches
       0: return -1.000000000000000;
       1: return -2.036650035073000;
       2: return -3.692974137304633;
       3: return -4.353162788050049;
       4: return -6.917614680418554;
       5: return -7.001372619757383;
       6: return -9.500983719365619;
       7: return -9.822964654887851;
       8: return -11.851583079120392;
       9: return -12.393321377282353;
      10: return -14.259426372933966;
      11: return -14.852920675443444;
      12: return -16.702718099601242;
      13: return -16.514466466800464;
      14: return -19.134794570592831;
      15: return -18.960789744323275;
      16: return -63.000000000000000;
      17: return -20.710057806027411;
      18: return -63.000000000000000;
      19: return -21.628249428489006;
      20: return -63.000000000000000;
      21: return -63.000000000000000;
      22: return -63.000000000000000;
      23: return -63.000000000000000;
      24: return -63.000000000000000;
      25: return -63.000000000000000;
      26: return -63.000000000000000;
      27: return -63.000000000000000;
      28: return -63.000000000000000;
      29: return -63.000000000000000;
      30: return -63.000000000000000;
      31: return -63.000000000000000;
      32: return -63.000000000000000;
      33: return -63.000000000000000;
      34: return -63.000000000000000;
      35: return -63.000000000000000;
      36: return -63.000000000000000;
      37: return -63.000000000000000;
      38: return -63.000000000000000;
      39: return -63.000000000000000;
      40: return -63.000000000000000;
      41: return -63.000000000000000;
      42: return -63.000000000000000;
      43: return -63.000000000000000;
      44: return -63.000000000000000;
      45: return -63.000000000000000;
      46: return -63.000000000000000;
      47: return -63.000000000000000;
      48: return -63.000000000000000;
      49: return -63.000000000000000;
      50: return -63.000000000000000;
      51: return -63.000000000000000;
      52: return -63.000000000000000;
      53: return -63.000000000000000;
      54: return -63.000000000000000;
      55: return -63.000000000000000;
      56: return -63.000000000000000;
      57: return -63.000000000000000;
      58: return -63.000000000000000;
      59: return -63.000000000000000;
      60: return -63.000000000000000;
      61: return -63.000000000000000;
      62: return -63.000000000000000;
      63: return -63.000000000000000;
      default: return -63;
   endcase
endfunction
