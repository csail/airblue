// generated by compute-ber.py
// table for rate 7 (exact)
// (computed without odd hints)

import Real::*;

function data_t get_ber_r7_log(Bit#(8) hint)
      provisos (RealLiteral#(data_t), Arith#(data_t));
   case (hint) matches
       0: return -1.000000000000000;
       1: return -1.191365780057514;
       2: return -1.410217776753495;
       3: return -1.630257465668733;
       4: return -1.934415522650261;
       5: return -2.169723228551087;
       6: return -2.582540357211471;
       7: return -2.813891820205739;
       8: return -3.383013421711915;
       9: return -3.581659171922587;
      10: return -4.318073409763133;
      11: return -4.436516305436519;
      12: return -5.380341360821678;
      13: return -5.382300236751637;
      14: return -6.533339357826147;
      15: return -6.345934966209284;
      16: return -7.745620476951301;
      17: return -7.332042008748800;
      18: return -8.997782012153092;
      19: return -8.380338705214584;
      20: return -10.280375394587217;
      21: return -9.409261451055253;
      22: return -11.521238087657329;
      23: return -10.779365923779086;
      24: return -12.735855341790680;
      25: return -11.676103999278238;
      26: return -14.060670627818800;
      27: return -12.609149874716230;
      28: return -15.135755797111877;
      29: return -13.634243841577469;
      30: return -15.733264568115786;
      31: return -63.000000000000000;
      32: return -17.264552557548473;
      33: return -63.000000000000000;
      34: return -63.000000000000000;
      35: return -63.000000000000000;
      36: return -63.000000000000000;
      37: return -63.000000000000000;
      38: return -63.000000000000000;
      39: return -63.000000000000000;
      40: return -63.000000000000000;
      41: return -63.000000000000000;
      42: return -63.000000000000000;
      43: return -63.000000000000000;
      44: return -63.000000000000000;
      45: return -63.000000000000000;
      46: return -63.000000000000000;
      47: return -63.000000000000000;
      48: return -63.000000000000000;
      49: return -63.000000000000000;
      50: return -63.000000000000000;
      51: return -63.000000000000000;
      52: return -63.000000000000000;
      53: return -63.000000000000000;
      54: return -63.000000000000000;
      55: return -63.000000000000000;
      56: return -63.000000000000000;
      57: return -63.000000000000000;
      58: return -63.000000000000000;
      59: return -63.000000000000000;
      60: return -63.000000000000000;
      61: return -63.000000000000000;
      62: return -63.000000000000000;
      63: return -63.000000000000000;
      default: return -63;
   endcase
endfunction
