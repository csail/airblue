// generated by compute-ber.py
// table for rate 1
// (computed without odd hints)

function BitErrorRate getBER_R1(SoftPhyHints hint);
   case (hint) matches
       0: return -1.0000000000;
       1: return -1.0000000000;
       2: return -1.2273409217;
       3: return -1.7042946352;
       4: return -2.2640590307;
       5: return -2.8884120609;
       6: return -3.5588309683;
       7: return -4.2600372214;
       8: return -4.9809311753;
       9: return -5.7140603783;
      10: return -6.4546585170;
      11: return -7.1997662284;
      12: return -7.9475786646;
      13: return -8.6970068521;
      14: return -9.4473979536;
      15: return -10.1983620901;
      16: return -10.9496669534;
      17: return -11.7011743105;
      18: return -12.4528019735;
      19: return -13.2045011002;
      20: return -13.9562426728;
      21: return -14.7080094548;
      22: return -15.4597912084;
      23: return -16.2115818534;
      24: return -16.9633777788;
      25: return -17.7151768399;
      26: return -18.4669777633;
      27: return -19.2187797926;
      28: return -19.9705824787;
      29: return -20.7223855548;
      30: return -21.4741888625;
      31: return -22.2259923078;
      32: return -22.9777958348;
      33: return -23.7295994103;
      34: return -24.4814030145;
      35: return -25.2332066359;
      36: return -25.9850102675;
      37: return -26.7368139051;
      38: return -27.4886175462;
      39: return -28.2404211895;
      40: return -28.9922248341;
      41: return -29.7440284794;
      42: return -30.4958321252;
      43: return -31.2476357712;
      44: return -31.9994394174;
      default: return -63;
   endcase
endfunction
