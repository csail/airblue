// generated by compute-ber.py
// table for rate 3 (exact)
// (computed without odd hints)

import Real::*;

function data_t get_ber_r3_log(Bit#(8) hint)
      provisos (RealLiteral#(data_t), Arith#(data_t));
   case (hint) matches
       0: return -1.000000000000000;
       1: return -1.812353834537644;
       2: return -2.963386716884308;
       3: return -3.896256285709370;
       4: return -5.524662941082885;
       5: return -6.270936607307813;
       6: return -8.150253602170402;
       7: return -8.607943218213931;
       8: return -10.735570684946309;
       9: return -10.863027513375410;
      10: return -13.872268841452433;
      11: return -13.172394788612525;
      12: return -16.501885133647420;
      13: return -15.416679904504369;
      14: return -19.740129904278177;
      15: return -17.327111212175655;
      16: return -23.325568493770010;
      17: return -19.687500286911963;
      18: return -28.111130335963672;
      19: return -21.251855097839389;
      20: return -63.000000000000000;
      21: return -63.000000000000000;
      22: return -63.000000000000000;
      23: return -63.000000000000000;
      24: return -63.000000000000000;
      25: return -63.000000000000000;
      26: return -63.000000000000000;
      27: return -63.000000000000000;
      28: return -63.000000000000000;
      29: return -63.000000000000000;
      30: return -63.000000000000000;
      31: return -63.000000000000000;
      32: return -63.000000000000000;
      33: return -63.000000000000000;
      34: return -63.000000000000000;
      35: return -63.000000000000000;
      36: return -63.000000000000000;
      37: return -63.000000000000000;
      38: return -63.000000000000000;
      39: return -63.000000000000000;
      40: return -63.000000000000000;
      41: return -63.000000000000000;
      42: return -63.000000000000000;
      43: return -63.000000000000000;
      44: return -63.000000000000000;
      45: return -63.000000000000000;
      46: return -63.000000000000000;
      47: return -63.000000000000000;
      48: return -63.000000000000000;
      49: return -63.000000000000000;
      50: return -63.000000000000000;
      51: return -63.000000000000000;
      52: return -63.000000000000000;
      53: return -63.000000000000000;
      54: return -63.000000000000000;
      55: return -63.000000000000000;
      56: return -63.000000000000000;
      57: return -63.000000000000000;
      58: return -63.000000000000000;
      59: return -63.000000000000000;
      60: return -63.000000000000000;
      61: return -63.000000000000000;
      62: return -63.000000000000000;
      63: return -63.000000000000000;
      default: return -63;
   endcase
endfunction
