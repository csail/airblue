// generated by compute-ber.py
// table for rate 7
// (computed without odd hints)

function BitErrorRate getBER_R7(SoftPhyHints hint);
   case (hint) matches
       0: return -1.0000000000;
       1: return -1.0000000000;
       2: return -1.0000000000;
       3: return -1.0000000000;
       4: return -1.0000000000;
       5: return -1.0446152951;
       6: return -1.3970082224;
       7: return -1.8117854641;
       8: return -2.2806732967;
       9: return -2.7931376060;
      10: return -3.3386377554;
      11: return -3.9080497617;
      12: return -4.4941938611;
      13: return -5.0917701477;
      14: return -5.6970305036;
      15: return -6.3073988515;
      16: return -6.9211378011;
      17: return -7.5370900898;
      18: return -8.1544911396;
      19: return -8.7728385004;
      20: return -9.3918031313;
      21: return -10.0111700415;
      22: return -10.6307989670;
      23: return -11.2505984852;
      24: return -11.8705090454;
      25: return -12.4904918732;
      26: return -13.1105217287;
      27: return -13.7305821852;
      28: return -14.3506625530;
      29: return -14.9707558760;
      30: return -15.5908576282;
      31: return -16.2109648648;
      32: return -16.8310756697;
      33: return -17.4511887962;
      34: return -18.0713034331;
      35: return -18.6914190528;
      36: return -19.3115353119;
      37: return -19.9316519870;
      38: return -20.5517689327;
      39: return -21.1718860546;
      40: return -21.7920032910;
      41: return -22.4121206020;
      42: return -23.0322379615;
      43: return -23.6523553525;
      44: return -24.2724727640;
      45: return -24.8925901889;
      46: return -25.5127076225;
      47: return -26.1328250618;
      48: return -26.7529425047;
      49: return -27.3730599500;
      50: return -27.9931773969;
      51: return -28.6132948448;
      52: return -29.2334122933;
      53: return -29.8535297423;
      54: return -30.4736471916;
      55: return -31.0937646410;
      56: return -31.7138820906;
      default: return -63;
   endcase
endfunction
