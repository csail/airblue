../../../parameters/WiFi/Macros.bsv