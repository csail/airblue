//----------------------------------------------------------------------//
// The MIT License 
// 
// Copyright (c) 2011 Kermin Fleming
// 
// Permission is hereby granted, free of charge, to any person 
// obtaining a copy of this software and associated documentation 
// files (the "Software"), to deal in the Software without 
// restriction, including without limitation the rights to use,
// copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the
// Software is furnished to do so, subject to the following conditions:
// 
// The above copyright notice and this permission notice shall be
// included in all copies or substantial portions of the Software.
// 
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
// EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES
// OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
// NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT
// HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY,
// WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
// FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR
// OTHER DEALINGS IN THE SOFTWARE.
//----------------------------------------------------------------------//

import FShow::*;
import Vector::*;

// This file contains airblue library-specific typeclasses
// and some general instances of these typeclasses

typeclass HasByteLength#(type a, numeric type m);
   function Bit#(m) byteLength(a value);
   function a setByteLength(a value, Bit#(m) length);
endtypeclass

instance HasByteLength#(Bit#(m), m);
   function Bit#(m) byteLength(Bit#(m) b) = b; 
   function Bit#(m) setByteLength(Bit#(m) b, Bit#(m) length);
      return length;
   endfunction
endinstance


typeclass EqualizerCtrl#(type a);
   function Bool initializeEqualizer(a value);
endtypeclass