// generated by compute-ber.py
// table for rate 6
// (computed without odd hints)

function BitErrorRate getBER_R6(SoftPhyHints hint);
   case (hint) matches
       0: return -1.0000000000;
       1: return -1.0000000000;
       2: return -1.0000000000;
       3: return -1.0000000000;
       4: return -1.0000000000;
       5: return -1.0000000000;
       6: return -1.1949412921;
       7: return -1.4915841185;
       8: return -1.8263684878;
       9: return -2.1949034521;
      10: return -2.5919468229;
      11: return -3.0121384357;
      12: return -3.4505297333;
      13: return -3.9028701496;
      14: return -4.3656942240;
      15: return -4.8362817465;
      16: return -5.3125555122;
      17: return -5.7929606473;
      18: return -6.2763498858;
      19: return -6.7618854245;
      20: return -7.2489599688;
      21: return -7.7371356412;
      22: return -8.2260979135;
      23: return -8.7156214703;
      24: return -9.2055452155;
      25: return -9.6957541270;
      26: return -10.1861661596;
      27: return -10.6767228315;
      28: return -11.1673824775;
      29: return -11.6581154238;
      30: return -12.1489005420;
      31: return -12.6397227914;
      32: return -13.1305714658;
      33: return -13.6214389452;
      34: return -14.1123198068;
      35: return -14.6032101912;
      36: return -15.0941073520;
      37: return -15.5850093348;
      38: return -16.0759147489;
      39: return -16.5668226046;
      40: return -17.0577321978;
      41: return -17.5486430273;
      42: return -18.0395547366;
      43: return -18.5304670718;
      44: return -19.0213798525;
      45: return -19.5122929502;
      46: return -20.0032062734;
      47: return -20.4941197570;
      48: return -20.9850333549;
      49: return -21.4759470341;
      50: return -21.9668607711;
      51: return -22.4577745492;
      52: return -22.9486883566;
      53: return -23.4396021849;
      54: return -23.9305160280;
      55: return -24.4214298816;
      56: return -24.9123437427;
      57: return -25.4032576092;
      58: return -25.8941714795;
      59: return -26.3850853524;
      60: return -26.8759992273;
      61: return -27.3669131036;
      62: return -27.8578269808;
      63: return -28.3487408588;
      64: return -28.8396547372;
      65: return -29.3305686160;
      66: return -29.8214824950;
      67: return -30.3123963742;
      68: return -30.8033102536;
      69: return -31.2942241330;
      70: return -31.7851380125;
      default: return -63;
   endcase
endfunction
