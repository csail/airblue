// generated by compute-ber.py
// table for rate 6 (exact)
// (computed without odd hints)

import Real::*;

function data_t get_ber_r6_log(Bit#(8) hint)
      provisos (RealLiteral#(data_t), Arith#(data_t));
   case (hint) matches
       0: return -1.001259510869769;
       1: return -1.132015740427657;
       2: return -1.282265914296657;
       3: return -1.421290686384904;
       4: return -1.625387718329333;
       5: return -1.774194750173572;
       6: return -2.042032508796354;
       7: return -2.203357512686926;
       8: return -2.557891396524304;
       9: return -2.723908757992830;
      10: return -3.180435268424036;
      11: return -3.346091348684866;
      12: return -3.914599835838715;
      13: return -4.071563682407961;
      14: return -4.749321458768335;
      15: return -4.851147345350777;
      16: return -5.660278394516863;
      17: return -5.716545224326494;
      18: return -6.627919349857358;
      19: return -6.608126037022275;
      20: return -7.641974785897178;
      21: return -7.449136070313407;
      22: return -8.675873805578355;
      23: return -8.412234132471530;
      24: return -9.752296654360478;
      25: return -9.490510959109827;
      26: return -10.791147389211238;
      27: return -10.303358874866134;
      28: return -11.916062251199893;
      29: return -11.468944530798634;
      30: return -13.020073998752903;
      31: return -12.007825427674247;
      32: return -14.301571682112746;
      33: return -14.968666793195208;
      34: return -16.003835860268794;
      35: return -63.000000000000000;
      36: return -16.405127956093480;
      37: return -63.000000000000000;
      38: return -18.890377101927072;
      39: return -63.000000000000000;
      40: return -63.000000000000000;
      41: return -63.000000000000000;
      42: return -63.000000000000000;
      43: return -63.000000000000000;
      44: return -63.000000000000000;
      45: return -63.000000000000000;
      46: return -63.000000000000000;
      47: return -63.000000000000000;
      48: return -63.000000000000000;
      49: return -63.000000000000000;
      50: return -63.000000000000000;
      51: return -63.000000000000000;
      52: return -63.000000000000000;
      53: return -63.000000000000000;
      54: return -63.000000000000000;
      55: return -63.000000000000000;
      56: return -63.000000000000000;
      57: return -63.000000000000000;
      58: return -63.000000000000000;
      59: return -63.000000000000000;
      60: return -63.000000000000000;
      61: return -63.000000000000000;
      62: return -63.000000000000000;
      63: return -63.000000000000000;
      default: return -63;
   endcase
endfunction
