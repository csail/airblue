********************************************************************
* Awb module specification
********************************************************************

%AWB_START

%name OFDM IFFT module
%desc OFDM IFFT module
%provides ofdm_ifft

%requires ofdm_fftifft

%attributes ofdm

%public IFFT.bsv

%AWB_END
 FParams.bsv FFTIFFT_Library.bsv