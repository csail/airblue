// generated by compute-ber.py
// table for rate 2
// (computed without odd hints)

function BitErrorRate getBER_R2(SoftPhyHints hint);
   case (hint) matches
       0: return -1.0000000000;
       1: return -1.3833831590;
       2: return -1.8460164051;
       3: return -2.3746102615;
       4: return -2.9545959698;
       5: return -3.5718628841;
       6: return -4.2147900470;
       7: return -4.8747438892;
       8: return -5.5457220107;
       9: return -6.2237248821;
      10: return -6.9061584327;
      11: return -7.5913685019;
      12: return -8.2783114462;
      13: return -8.9663331683;
      14: return -9.6550254082;
      15: return -10.3441340010;
      16: return -11.0335009671;
      17: return -11.7230282096;
      18: return -12.4126548527;
      19: return -13.1023431333;
      20: return -13.7920696314;
      21: return -14.4818198244;
      22: return -15.1715847077;
      23: return -15.8613586986;
      24: return -16.5511383357;
      25: return -17.2409214733;
      26: return -17.9307067809;
      27: return -18.6204934340;
      28: return -19.3102809210;
      29: return -20.0000689251;
      30: return -20.6898572498;
      31: return -21.3796457731;
      32: return -22.0694344197;
      33: return -22.7592231427;
      34: return -23.4490119130;
      35: return -24.1388007126;
      36: return -24.8285895305;
      37: return -25.5183783596;
      38: return -26.2081671957;
      39: return -26.8979560362;
      40: return -27.5877448793;
      41: return -28.2775337241;
      42: return -28.9673225700;
      43: return -29.6571114165;
      44: return -30.3469002634;
      45: return -31.0366891105;
      46: return -31.7264779578;
      default: return -63;
   endcase
endfunction
