// generated by compute-ber.py
// table for rate 2 (exact)
// (computed without odd hints)

import Real::*;

function data_t get_ber_r2_log(Bit#(8) hint)
      provisos (RealLiteral#(data_t), Arith#(data_t));
   case (hint) matches
       0: return -1.000000000000000;
       1: return -1.904671795811353;
       2: return -3.790730753718377;
       3: return -4.902210315620936;
       4: return -7.524782537484684;
       5: return -7.816047061659566;
       6: return -11.734370919662975;
       7: return -11.528161048833141;
       8: return -15.162902664709245;
       9: return -13.758847803108321;
      10: return -63.000000000000000;
      11: return -16.666404328413176;
      12: return -63.000000000000000;
      13: return -63.000000000000000;
      14: return -63.000000000000000;
      15: return -63.000000000000000;
      16: return -63.000000000000000;
      17: return -63.000000000000000;
      18: return -63.000000000000000;
      19: return -63.000000000000000;
      20: return -63.000000000000000;
      21: return -63.000000000000000;
      22: return -63.000000000000000;
      23: return -63.000000000000000;
      24: return -63.000000000000000;
      25: return -63.000000000000000;
      26: return -63.000000000000000;
      27: return -63.000000000000000;
      28: return -63.000000000000000;
      29: return -63.000000000000000;
      30: return -63.000000000000000;
      31: return -63.000000000000000;
      32: return -63.000000000000000;
      33: return -63.000000000000000;
      34: return -63.000000000000000;
      35: return -63.000000000000000;
      36: return -63.000000000000000;
      37: return -63.000000000000000;
      38: return -63.000000000000000;
      39: return -63.000000000000000;
      40: return -63.000000000000000;
      41: return -63.000000000000000;
      42: return -63.000000000000000;
      43: return -63.000000000000000;
      44: return -63.000000000000000;
      45: return -63.000000000000000;
      46: return -63.000000000000000;
      47: return -63.000000000000000;
      48: return -63.000000000000000;
      49: return -63.000000000000000;
      50: return -63.000000000000000;
      51: return -63.000000000000000;
      52: return -63.000000000000000;
      53: return -63.000000000000000;
      54: return -63.000000000000000;
      55: return -63.000000000000000;
      56: return -63.000000000000000;
      57: return -63.000000000000000;
      58: return -63.000000000000000;
      59: return -63.000000000000000;
      60: return -63.000000000000000;
      61: return -63.000000000000000;
      62: return -63.000000000000000;
      63: return -63.000000000000000;
      default: return -63;
   endcase
endfunction
