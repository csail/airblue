// generated by compute-ber.py
// table for rate 4
// (computed without odd hints)

function BitErrorRate getBER_R4(SoftPhyHints hint);
   case (hint) matches
       0: return -1.0000000000;
       1: return -1.0000000000;
       2: return -1.0000000000;
       3: return -1.0000000000;
       4: return -1.0000000000;
       5: return -1.1973395887;
       6: return -1.4449196396;
       7: return -1.7199784506;
       8: return -2.0200560518;
       9: return -2.3421404008;
      10: return -2.6830018583;
      11: return -3.0394727473;
      12: return -3.4086408659;
      13: return -3.7879558447;
      14: return -4.1752652133;
      15: return -4.5688028540;
      16: return -4.9671505228;
      17: return -5.3691878556;
      18: return -5.7740407662;
      19: return -6.1810337233;
      20: return -6.5896483662;
      21: return -6.9994890797;
      22: return -7.4102551553;
      23: return -7.8217187240;
      24: return -8.2337075109;
      25: return -8.6460914979;
      26: return -9.0587726869;
      27: return -9.4716772863;
      28: return -9.8847497733;
      29: return -10.2979483935;
      30: return -10.7112417604;
      31: return -11.1246062879;
      32: return -11.5380242561;
      33: return -11.9514823545;
      34: return -12.3649705861;
      35: return -12.7784814434;
      36: return -13.1920092888;
      37: return -13.6055498890;
      38: return -14.0191000656;
      39: return -14.4326574320;
      40: return -14.8462201964;
      41: return -15.2597870134;
      42: return -15.6733568731;
      43: return -16.0869290171;
      44: return -16.5005028761;
      45: return -16.9140780226;
      46: return -17.3276541358;
      47: return -17.7412309747;
      48: return -18.1548083584;
      49: return -18.5683861512;
      50: return -18.9819642510;
      51: return -19.3955425815;
      52: return -19.8091210850;
      53: return -20.2226997184;
      54: return -20.6362784495;
      55: return -21.0498572537;
      56: return -21.4634361130;
      57: return -21.8770150135;
      58: return -22.2905939451;
      59: return -22.7041728999;
      60: return -23.1177518722;
      61: return -23.5313308575;
      62: return -23.9449098528;
      63: return -24.3584888554;
      64: return -24.7720678636;
      65: return -25.1856468759;
      66: return -25.5992258914;
      67: return -26.0128049092;
      68: return -26.4263839288;
      69: return -26.8399629497;
      70: return -27.2535419716;
      71: return -27.6671209943;
      72: return -28.0807000175;
      73: return -28.4942790411;
      74: return -28.9078580651;
      75: return -29.3214370892;
      76: return -29.7350161136;
      77: return -30.1485951381;
      78: return -30.5621741627;
      79: return -30.9757531873;
      80: return -31.3893322121;
      81: return -31.8029112368;
      default: return -63;
   endcase
endfunction
