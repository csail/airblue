// generated by compute-ber.py
// table for rate 5
// (computed without odd hints)

function BitErrorRate getBER_R5(SoftPhyHints hint);
   case (hint) matches
       0: return -1.0000000000;
       1: return -1.0000000000;
       2: return -1.0000000000;
       3: return -1.0000000000;
       4: return -1.0000000000;
       5: return -1.3050564991;
       6: return -1.7390982912;
       7: return -2.2378736135;
       8: return -2.7884216577;
       9: return -3.3775122323;
      10: return -3.9937852918;
      11: return -4.6285031901;
      12: return -5.2754104306;
      13: return -5.9302326153;
      14: return -6.5901356102;
      15: return -7.2532761053;
      16: return -7.9184698332;
      17: return -8.5849618333;
      18: return -9.2522731847;
      19: return -9.9201010176;
      20: return -10.5882541710;
      21: return -11.2566121394;
      22: return -11.9250990165;
      23: return -12.5936670123;
      24: return -13.2622860476;
      25: return -13.9309371945;
      26: return -14.5996085436;
      27: return -15.2682926018;
      28: return -15.9369846552;
      29: return -16.6056817383;
      30: return -17.2743819854;
      31: return -17.9430842230;
      32: return -18.6117877127;
      33: return -19.2804919901;
      34: return -19.9491967630;
      35: return -20.6179018476;
      36: return -21.2866071283;
      37: return -21.9553125323;
      38: return -22.6240180139;
      39: return -23.2927235444;
      40: return -23.9614291056;
      41: return -24.6301346860;
      42: return -25.2988402787;
      43: return -25.9675458789;
      44: return -26.6362514840;
      45: return -27.3049570921;
      46: return -27.9736627021;
      47: return -28.6423683133;
      48: return -29.3110739253;
      49: return -29.9797795377;
      50: return -30.6484851505;
      51: return -31.3171907634;
      52: return -31.9858963764;
      default: return -63;
   endcase
endfunction
