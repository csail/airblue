
typedef 32 FFTIFFTSz;

typedef 4  TXFPFPrec;
typedef 14  TXFPIPrec;