// generated by compute-ber.py
// table for rate 3
// (computed without odd hints)

function BitErrorRate getBER_R3(SoftPhyHints hint);
   case (hint) matches
       0: return -1.0000000000;
       1: return -1.0000000000;
       2: return -1.0000000000;
       3: return -1.4110583859;
       4: return -1.9475802975;
       5: return -2.5656164005;
       6: return -3.2436893980;
       7: return -3.9624191106;
       8: return -4.7071295954;
       9: return -5.4678290304;
      10: return -6.2381404975;
      11: return -7.0141490405;
      12: return -7.7935058709;
      13: return -8.5748207937;
      14: return -9.3572774859;
      15: return -10.1403988157;
      16: return -10.9239066564;
      17: return -11.7076391375;
      18: return -12.4915021361;
      19: return -13.2754409515;
      20: return -14.0594238034;
      21: return -14.8434322312;
      22: return -15.6274555126;
      23: return -16.4114874204;
      24: return -17.1955243380;
      25: return -17.9795641648;
      26: return -18.7636056813;
      27: return -19.5476481789;
      28: return -20.3316912464;
      29: return -21.1157346448;
      30: return -21.8997782354;
      31: return -22.6838219375;
      32: return -23.4678657045;
      33: return -24.2519095091;
      34: return -25.0359533356;
      35: return -25.8199971748;
      36: return -26.6040410213;
      37: return -27.3880848722;
      38: return -28.1721287255;
      39: return -28.9561725802;
      40: return -29.7402164358;
      41: return -30.5242602919;
      42: return -31.3083041483;
      default: return -63;
   endcase
endfunction
