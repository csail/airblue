import DataTypes::*;
import Controls::*;
import Interfaces::*;
import Typeclasses::*;
export DataTypes::*;
export Controls::*;
export Interfaces::*;
export Typeclasses::*;

