// bsv libraries
import Vector::*;
import FIFO::*;
import Connectable::*;

// portz libraries
import CtrlMux::*;
import Portal::*;
import Leds::*;
import MemTypes::*;
import MemPortal::*;

// defined by user
import ScramblerTest::*;

// generated by tool
import ScramblerIndicationProxy::*;
import ScramblerRequestWrapper::*;

module mkConnectalTop(StdConnectalTop#(PhysAddrWidth));

   // instantiate user portals
   ScramblerIndicationProxy scramblerIndicationProxy <- mkScramblerIndicationProxy(ScramblerIndicationPortal);
   ScramblerRequest scramblerTest <- mkScramblerTest(scramblerIndicationProxy.ifc);
   ScramblerRequestWrapper scramblerRequestWrapper <- mkScramblerRequestWrapper(ScramblerRequestPortal,scramblerTest);
   
   Vector#(2,StdPortal) portals;
   portals[0] = scramblerRequestWrapper.portalIfc;
   portals[1] = scramblerIndicationProxy.portalIfc;

   // instantiate system directory
   let ctrl_mux <- mkSlaveMux(portals);
   
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = nil;
   interface leds = default_leds;

endmodule : mkConnectalTop


