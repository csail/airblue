../../Viterbi/src/Macros.bsv