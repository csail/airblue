//This file contains architecture parameters relevant to the FFT

typedef 4             FFTIFFTNoBfly;

