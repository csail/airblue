../../common/src/Macros.bsv