import Vector::*;

import ofdm_base::*;

//
// import EHRReg::*;
/////////////////////////////////////////////////////////////
// Interface
// Name: StreamFIFO
// Ptrs: sz, s_sz, data_t
// Dscr: A fifo that can enq and deq arbitrary no. of 
//       elements
/////////////////////////////////////////////////////////////
interface StreamFIFO#(numeric type sz,     // buffer sz
		      numeric type s_sz,   // shift sz
		      type data_t);        // basic data unit
      method Action enq(Bit#(s_sz) i_s_sz, 
			Vector#(sz, data_t) i_msg);
      method Vector#(sz, data_t) first();
      method Action deq(Bit#(s_sz) o_s_sz); 
      method Action clear();
      method Bool notEmpty(Bit#(s_sz) o_s_sz); // canDeq?
      method Bool notFull(Bit#(s_sz) i_s_sz);  // canEnq?
      method Bit#(s_sz) usage(); // no of slots used
      method Bit#(s_sz) free(); // no of slots unused
endinterface

//////////////////////////////////////////////////////////////
// Functions
/////////////////////////////////////////////////////////////
// shift towards higher index
function Vector#(sz,data_t) shiftLeftBy(Vector#(sz,data_t) inVec,
					Bit#(s_sz) shiftBy)
   provisos (Add#(sz,1,szp1),
	     Log#(szp1,s_sz),
	     Bits#(data_t,data_sz));
   
   function Vector#(sz,data_t) stageFunc(Vector#(sz,data_t) iVec,
					 Tuple2#(Bit#(1),Nat) ctrl);
      return (tpl_1(ctrl) == 1) ? 
             unpack(pack(iVec) << tpl_2(ctrl)) : 
             iVec;
   endfunction
   
   Nat dataSz = fromInteger(valueOf(data_sz));
   Vector#(s_sz,Bit#(1)) shiftVec = unpack(shiftBy);
   Vector#(s_sz,Nat) natVec0 = genWith(fromInteger);
   Vector#(s_sz,Nat) natVec1 = map(\<< (1),natVec0);
   Vector#(s_sz,Nat) natVec2 = map(\* (dataSz),natVec1);
   let ctrlVec = zip(shiftVec, natVec2);
   return foldl(stageFunc,inVec,ctrlVec);
   
endfunction

// shift towards lower index
function Vector#(sz,data_t) shiftRightBy(Vector#(sz,data_t) inVec,
					 Bit#(s_sz) shiftBy)
   provisos (Add#(sz,1,szp1),
	     Log#(szp1,s_sz),
	     Bits#(data_t,data_sz));
   
   function Vector#(sz,data_t) stageFunc(Vector#(sz,data_t) iVec,
					 Tuple2#(Bit#(1),Nat) ctrl);
      return (tpl_1(ctrl) == 1) ? 
             unpack(pack(iVec) >> tpl_2(ctrl)) : 
             iVec;
   endfunction
   
   Nat dataSz = fromInteger(valueOf(data_sz));
   Vector#(s_sz,Bit#(1)) shiftVec = unpack(shiftBy);
   Vector#(s_sz,Nat) natVec0 = genWith(fromInteger);
   Vector#(s_sz,Nat) natVec1 = map(\<< (1),natVec0);
   Vector#(s_sz,Nat) natVec2 = map(\* (dataSz),natVec1);
   let ctrlVec = zip(shiftVec, natVec2);
   return foldl(stageFunc,inVec,ctrlVec);
   
endfunction


////////////////////////////////////////////////////////////////////
// Module
// Name: mkStreamFIFO
// Ptrs: 
// Dscr: Create an instance of StreamFIFO which is implemented with
//       shifting approach
// Notes: To enq/deq, caller needs to check notFull/notEmpty 
//        explicitly  
///////////////////////////////////////////////////////////////////
module mkStreamFIFO(StreamFIFO#(sz, s_sz, data_t))
   provisos (Add#(sz,1,szp1),
	     Log#(szp1,s_sz),
	     Bits#(data_t,data_sz));
   
   Bit#(s_sz) maxTail = fromInteger(valueOf(sz));
   EHRReg#(2,Vector#(sz,data_t)) buffer <- mkEHRReg(newVector);       
   EHRReg#(2,Bit#(s_sz)) tail <- mkEHRReg(0); // equal to usage
   
   function data_t selTuple(Tuple3#(Bool,data_t,data_t) tup);
      return tpl_1(tup) ? tpl_2(tup) : tpl_3(tup);
   endfunction

   method Action enq(Bit#(s_sz) i_s_sz, 
		     Vector#(sz, data_t) i_msg);
      let buffer0 = buffer[1];
      let buffer1 = shiftLeftBy(i_msg, tail[1]);
      Vector#(sz, Bit#(s_sz)) idxVec = genWith(fromInteger);
      Vector#(sz, Bool) selBuffer = map(\> (tail[1]), idxVec);
      let zipBuffer = zip3(selBuffer,buffer0,buffer1);
      let newBuffer = map(selTuple,zipBuffer);
      buffer[1] <= newBuffer;
      tail[1] <= tail[1] + i_s_sz;
   endmethod
   
   method Vector#(sz, data_t) first(); 
      return buffer[0];
   endmethod
   
   method Action deq(Bit#(s_sz) o_s_sz);
      buffer[0] <= shiftRightBy(buffer[0], o_s_sz);
      tail[0] <= tail[0] - o_s_sz;
   endmethod
   
   method Action clear();
      tail[1] <= 0;
   endmethod
   
   method Bool notEmpty(Bit#(s_sz) o_s_sz);
      return tail[0] >= o_s_sz;
   endmethod
   
   method Bool notFull(Bit#(s_sz) i_s_sz);
      return tail[0] <= maxTail - i_s_sz;
   endmethod
   
   method Bit#(s_sz) usage();
      return tail[0];
   endmethod
   
   method Bit#(s_sz) free();
      return maxTail - tail[0];
   endmethod
endmodule

////////////////////////////////////////////////////////////////////
// Module
// Name: mkStreamLFIFO
// Ptrs: 
// Dscr: Create an instance of StreamFIFO which is implemented with
//       shifting approach, can deq and enq parallelly when it is full
// Notes: To enq/deq, caller needs to check notFull/notEmpty 
//        explicitly  
///////////////////////////////////////////////////////////////////
module mkStreamLFIFO(StreamFIFO#(sz, s_sz, data_t))
   provisos (Add#(sz,1,szp1),
	     Log#(szp1,s_sz),
	     Bits#(data_t,data_sz));
   
   Bit#(s_sz) maxTail = fromInteger(valueOf(sz));
   EHRReg#(2,Vector#(sz,data_t)) buffer <- mkEHRReg(newVector);       
   EHRReg#(2,Bit#(s_sz)) tail <- mkEHRReg(0); // equal to usage
   
   function data_t selTuple(Tuple3#(Bool,data_t,data_t) tup);
      return tpl_1(tup) ? tpl_2(tup) : tpl_3(tup);
   endfunction

   method Action enq(Bit#(s_sz) i_s_sz, 
		     Vector#(sz, data_t) i_msg);
      let buffer0 = buffer[1];
      let buffer1 = shiftLeftBy(i_msg, tail[1]);
      Vector#(sz, Bit#(s_sz)) idxVec = genWith(fromInteger);
      Vector#(sz, Bool) selBuffer = map(\> (tail[1]), idxVec);
      let zipBuffer = zip3(selBuffer,buffer0,buffer1);
      let newBuffer = map(selTuple,zipBuffer);
      buffer[1] <= newBuffer;
      tail[1] <= tail[1] + i_s_sz;
   endmethod
   
   method Vector#(sz, data_t) first(); 
      return buffer[0];
   endmethod
   
   method Action deq(Bit#(s_sz) o_s_sz);
      buffer[0] <= shiftRightBy(buffer[0], o_s_sz);
      tail[0] <= tail[0] - o_s_sz;
   endmethod
   
   method Action clear();
      tail[1] <= 0;
   endmethod
   
   method Bool notEmpty(Bit#(s_sz) o_s_sz);
      return tail[0] >= o_s_sz;
   endmethod
   
   method Bool notFull(Bit#(s_sz) i_s_sz);
      return tail[1] <= maxTail - i_s_sz; // slower ready signal 
   endmethod

   method Bit#(s_sz) usage();
      return tail[0];
   endmethod
   
   method Bit#(s_sz) free();
      return maxTail - tail[1];
   endmethod   
endmodule

