import Vector::*;

function fxptType getScale(Bit#(12) scale)
provisos(RealLiteral#(fxptType));
Vector#(4096,fxptType) scaleFactors = newVector;
scaleFactors[4095] = 0.0;
scaleFactors[4094] = 0.0;
scaleFactors[4093] = 0.0;
scaleFactors[4092] = 0.0;
scaleFactors[4091] = 0.0;
scaleFactors[4090] = 0.0;
scaleFactors[4089] = 0.0;
scaleFactors[4088] = 0.0;
scaleFactors[4087] = 0.0;
scaleFactors[4086] = 0.0;
scaleFactors[4085] = 0.0;
scaleFactors[4084] = 0.0;
scaleFactors[4083] = 0.0;
scaleFactors[4082] = 0.0;
scaleFactors[4081] = 0.0;
scaleFactors[4080] = 0.0;
scaleFactors[4079] = 0.0;
scaleFactors[4078] = 0.0;
scaleFactors[4077] = 0.0;
scaleFactors[4076] = 0.0;
scaleFactors[4075] = 0.0;
scaleFactors[4074] = 0.0;
scaleFactors[4073] = 0.0;
scaleFactors[4072] = 0.0;
scaleFactors[4071] = 0.0;
scaleFactors[4070] = 0.0;
scaleFactors[4069] = 0.0;
scaleFactors[4068] = 0.0;
scaleFactors[4067] = 0.0;
scaleFactors[4066] = 0.0;
scaleFactors[4065] = 0.0;
scaleFactors[4064] = 0.0;
scaleFactors[4063] = 0.0;
scaleFactors[4062] = 0.0;
scaleFactors[4061] = 0.0;
scaleFactors[4060] = 0.0;
scaleFactors[4059] = 0.0;
scaleFactors[4058] = 0.0;
scaleFactors[4057] = 0.0;
scaleFactors[4056] = 0.0;
scaleFactors[4055] = 0.0;
scaleFactors[4054] = 0.0;
scaleFactors[4053] = 0.0;
scaleFactors[4052] = 0.0;
scaleFactors[4051] = 0.0;
scaleFactors[4050] = 0.0;
scaleFactors[4049] = 0.0;
scaleFactors[4048] = 0.0;
scaleFactors[4047] = 0.0;
scaleFactors[4046] = 0.0;
scaleFactors[4045] = 0.0;
scaleFactors[4044] = 0.0;
scaleFactors[4043] = 0.0;
scaleFactors[4042] = 0.0;
scaleFactors[4041] = 0.0;
scaleFactors[4040] = 0.0;
scaleFactors[4039] = 0.0;
scaleFactors[4038] = 0.0;
scaleFactors[4037] = 0.0;
scaleFactors[4036] = 0.0;
scaleFactors[4035] = 0.0;
scaleFactors[4034] = 0.0;
scaleFactors[4033] = 0.0;
scaleFactors[4032] = 0.0;
scaleFactors[4031] = 0.0;
scaleFactors[4030] = 0.0;
scaleFactors[4029] = 0.0;
scaleFactors[4028] = 0.0;
scaleFactors[4027] = 0.0;
scaleFactors[4026] = 0.0;
scaleFactors[4025] = 0.0;
scaleFactors[4024] = 0.0;
scaleFactors[4023] = 0.0;
scaleFactors[4022] = 0.0;
scaleFactors[4021] = 0.0;
scaleFactors[4020] = 0.0;
scaleFactors[4019] = 0.0;
scaleFactors[4018] = 0.0;
scaleFactors[4017] = 0.0;
scaleFactors[4016] = 0.0;
scaleFactors[4015] = 0.0;
scaleFactors[4014] = 0.0;
scaleFactors[4013] = 0.0;
scaleFactors[4012] = 0.0;
scaleFactors[4011] = 0.0;
scaleFactors[4010] = 0.0;
scaleFactors[4009] = 0.0;
scaleFactors[4008] = 0.0;
scaleFactors[4007] = 0.0;
scaleFactors[4006] = 0.0;
scaleFactors[4005] = 0.0;
scaleFactors[4004] = 0.0;
scaleFactors[4003] = 0.0;
scaleFactors[4002] = 0.0;
scaleFactors[4001] = 0.0;
scaleFactors[4000] = 0.0;
scaleFactors[3999] = 0.0;
scaleFactors[3998] = 0.0;
scaleFactors[3997] = 0.0;
scaleFactors[3996] = 0.0;
scaleFactors[3995] = 0.0;
scaleFactors[3994] = 0.0;
scaleFactors[3993] = 0.0;
scaleFactors[3992] = 0.0;
scaleFactors[3991] = 0.0;
scaleFactors[3990] = 0.0;
scaleFactors[3989] = 0.0;
scaleFactors[3988] = 0.0;
scaleFactors[3987] = 0.0;
scaleFactors[3986] = 0.0;
scaleFactors[3985] = 0.0;
scaleFactors[3984] = 0.0;
scaleFactors[3983] = 0.0;
scaleFactors[3982] = 0.0;
scaleFactors[3981] = 0.0;
scaleFactors[3980] = 0.0;
scaleFactors[3979] = 0.0;
scaleFactors[3978] = 0.0;
scaleFactors[3977] = 0.0;
scaleFactors[3976] = 0.0;
scaleFactors[3975] = 0.0;
scaleFactors[3974] = 0.0;
scaleFactors[3973] = 0.0;
scaleFactors[3972] = 0.0;
scaleFactors[3971] = 0.0;
scaleFactors[3970] = 0.0;
scaleFactors[3969] = 0.0;
scaleFactors[3968] = 0.0;
scaleFactors[3967] = 0.0;
scaleFactors[3966] = 0.0;
scaleFactors[3965] = 0.0;
scaleFactors[3964] = 0.0;
scaleFactors[3963] = 0.0;
scaleFactors[3962] = 0.0;
scaleFactors[3961] = 0.0;
scaleFactors[3960] = 0.0;
scaleFactors[3959] = 0.0;
scaleFactors[3958] = 0.0;
scaleFactors[3957] = 0.0;
scaleFactors[3956] = 0.0;
scaleFactors[3955] = 0.0;
scaleFactors[3954] = 0.0;
scaleFactors[3953] = 0.0;
scaleFactors[3952] = 0.0;
scaleFactors[3951] = 0.0;
scaleFactors[3950] = 0.0;
scaleFactors[3949] = 0.0;
scaleFactors[3948] = 0.0;
scaleFactors[3947] = 0.0;
scaleFactors[3946] = 0.0;
scaleFactors[3945] = 0.0;
scaleFactors[3944] = 0.0;
scaleFactors[3943] = 0.0;
scaleFactors[3942] = 0.0;
scaleFactors[3941] = 0.0;
scaleFactors[3940] = 0.0;
scaleFactors[3939] = 0.0;
scaleFactors[3938] = 0.0;
scaleFactors[3937] = 0.0;
scaleFactors[3936] = 0.0;
scaleFactors[3935] = 0.0;
scaleFactors[3934] = 0.0;
scaleFactors[3933] = 0.0;
scaleFactors[3932] = 0.0;
scaleFactors[3931] = 0.0;
scaleFactors[3930] = 0.0;
scaleFactors[3929] = 0.0;
scaleFactors[3928] = 0.0;
scaleFactors[3927] = 0.0;
scaleFactors[3926] = 0.0;
scaleFactors[3925] = 0.0;
scaleFactors[3924] = 0.0;
scaleFactors[3923] = 0.0;
scaleFactors[3922] = 0.0;
scaleFactors[3921] = 0.0;
scaleFactors[3920] = 0.0;
scaleFactors[3919] = 0.0;
scaleFactors[3918] = 0.0;
scaleFactors[3917] = 0.0;
scaleFactors[3916] = 0.0;
scaleFactors[3915] = 0.0;
scaleFactors[3914] = 0.0;
scaleFactors[3913] = 0.0;
scaleFactors[3912] = 0.0;
scaleFactors[3911] = 0.0;
scaleFactors[3910] = 0.0;
scaleFactors[3909] = 0.0;
scaleFactors[3908] = 0.0;
scaleFactors[3907] = 0.0;
scaleFactors[3906] = 0.0;
scaleFactors[3905] = 0.0;
scaleFactors[3904] = 0.0;
scaleFactors[3903] = 0.0;
scaleFactors[3902] = 0.0;
scaleFactors[3901] = 0.0;
scaleFactors[3900] = 0.0;
scaleFactors[3899] = 0.0;
scaleFactors[3898] = 0.0;
scaleFactors[3897] = 0.0;
scaleFactors[3896] = 0.0;
scaleFactors[3895] = 0.0;
scaleFactors[3894] = 0.0;
scaleFactors[3893] = 0.0;
scaleFactors[3892] = 0.0;
scaleFactors[3891] = 0.0;
scaleFactors[3890] = 0.0;
scaleFactors[3889] = 0.0;
scaleFactors[3888] = 0.0;
scaleFactors[3887] = 0.0;
scaleFactors[3886] = 0.0;
scaleFactors[3885] = 0.0;
scaleFactors[3884] = 0.0;
scaleFactors[3883] = 0.0;
scaleFactors[3882] = 0.0;
scaleFactors[3881] = 0.0;
scaleFactors[3880] = 0.0;
scaleFactors[3879] = 0.0;
scaleFactors[3878] = 0.0;
scaleFactors[3877] = 0.0;
scaleFactors[3876] = 0.0;
scaleFactors[3875] = 0.0;
scaleFactors[3874] = 0.0;
scaleFactors[3873] = 0.0;
scaleFactors[3872] = 0.0;
scaleFactors[3871] = 0.0;
scaleFactors[3870] = 0.0;
scaleFactors[3869] = 0.0;
scaleFactors[3868] = 0.0;
scaleFactors[3867] = 0.0;
scaleFactors[3866] = 0.0;
scaleFactors[3865] = 0.0;
scaleFactors[3864] = 0.0;
scaleFactors[3863] = 0.0;
scaleFactors[3862] = 0.0;
scaleFactors[3861] = 0.0;
scaleFactors[3860] = 0.0;
scaleFactors[3859] = 0.0;
scaleFactors[3858] = 0.0;
scaleFactors[3857] = 0.0;
scaleFactors[3856] = 0.0;
scaleFactors[3855] = 0.0;
scaleFactors[3854] = 0.0;
scaleFactors[3853] = 0.0;
scaleFactors[3852] = 0.0;
scaleFactors[3851] = 0.0;
scaleFactors[3850] = 0.0;
scaleFactors[3849] = 0.0;
scaleFactors[3848] = 0.0;
scaleFactors[3847] = 0.0;
scaleFactors[3846] = 0.0;
scaleFactors[3845] = 0.0;
scaleFactors[3844] = 0.0;
scaleFactors[3843] = 0.0;
scaleFactors[3842] = 0.0;
scaleFactors[3841] = 0.0;
scaleFactors[3840] = 0.0;
scaleFactors[3839] = 0.0;
scaleFactors[3838] = 0.0;
scaleFactors[3837] = 0.0;
scaleFactors[3836] = 0.0;
scaleFactors[3835] = 0.0;
scaleFactors[3834] = 0.0;
scaleFactors[3833] = 0.0;
scaleFactors[3832] = 0.0;
scaleFactors[3831] = 0.0;
scaleFactors[3830] = 0.0;
scaleFactors[3829] = 0.0;
scaleFactors[3828] = 0.0;
scaleFactors[3827] = 0.0;
scaleFactors[3826] = 0.0;
scaleFactors[3825] = 0.0;
scaleFactors[3824] = 0.0;
scaleFactors[3823] = 0.0;
scaleFactors[3822] = 0.0;
scaleFactors[3821] = 0.0;
scaleFactors[3820] = 0.0;
scaleFactors[3819] = 0.0;
scaleFactors[3818] = 0.0;
scaleFactors[3817] = 0.0;
scaleFactors[3816] = 0.0;
scaleFactors[3815] = 0.0;
scaleFactors[3814] = 0.0;
scaleFactors[3813] = 0.0;
scaleFactors[3812] = 0.0;
scaleFactors[3811] = 0.0;
scaleFactors[3810] = 0.0;
scaleFactors[3809] = 0.0;
scaleFactors[3808] = 0.0;
scaleFactors[3807] = 0.0;
scaleFactors[3806] = 0.0;
scaleFactors[3805] = 0.0;
scaleFactors[3804] = 0.0;
scaleFactors[3803] = 0.0;
scaleFactors[3802] = 0.0;
scaleFactors[3801] = 0.0;
scaleFactors[3800] = 0.0;
scaleFactors[3799] = 0.0;
scaleFactors[3798] = 0.0;
scaleFactors[3797] = 0.0;
scaleFactors[3796] = 0.0;
scaleFactors[3795] = 0.0;
scaleFactors[3794] = 0.0;
scaleFactors[3793] = 0.0;
scaleFactors[3792] = 0.0;
scaleFactors[3791] = 0.0;
scaleFactors[3790] = 0.0;
scaleFactors[3789] = 0.0;
scaleFactors[3788] = 0.0;
scaleFactors[3787] = 0.0;
scaleFactors[3786] = 0.0;
scaleFactors[3785] = 0.0;
scaleFactors[3784] = 0.0;
scaleFactors[3783] = 0.0;
scaleFactors[3782] = 0.0;
scaleFactors[3781] = 0.0;
scaleFactors[3780] = 0.0;
scaleFactors[3779] = 0.0;
scaleFactors[3778] = 0.0;
scaleFactors[3777] = 0.0;
scaleFactors[3776] = 0.0;
scaleFactors[3775] = 0.0;
scaleFactors[3774] = 0.0;
scaleFactors[3773] = 0.0;
scaleFactors[3772] = 0.0;
scaleFactors[3771] = 0.0;
scaleFactors[3770] = 0.0;
scaleFactors[3769] = 0.0;
scaleFactors[3768] = 0.0;
scaleFactors[3767] = 0.0;
scaleFactors[3766] = 0.0;
scaleFactors[3765] = 0.0;
scaleFactors[3764] = 0.0;
scaleFactors[3763] = 0.0;
scaleFactors[3762] = 0.0;
scaleFactors[3761] = 0.0;
scaleFactors[3760] = 0.0;
scaleFactors[3759] = 0.0;
scaleFactors[3758] = 0.0;
scaleFactors[3757] = 0.0;
scaleFactors[3756] = 0.0;
scaleFactors[3755] = 0.0;
scaleFactors[3754] = 0.0;
scaleFactors[3753] = 0.0;
scaleFactors[3752] = 0.0;
scaleFactors[3751] = 0.0;
scaleFactors[3750] = 0.0;
scaleFactors[3749] = 0.0;
scaleFactors[3748] = 0.0;
scaleFactors[3747] = 0.0;
scaleFactors[3746] = 0.0;
scaleFactors[3745] = 0.0;
scaleFactors[3744] = 0.0;
scaleFactors[3743] = 0.0;
scaleFactors[3742] = 0.0;
scaleFactors[3741] = 0.0;
scaleFactors[3740] = 0.0;
scaleFactors[3739] = 0.0;
scaleFactors[3738] = 0.0;
scaleFactors[3737] = 0.0;
scaleFactors[3736] = 0.0;
scaleFactors[3735] = 0.0;
scaleFactors[3734] = 0.0;
scaleFactors[3733] = 0.0;
scaleFactors[3732] = 0.0;
scaleFactors[3731] = 0.0;
scaleFactors[3730] = 0.0;
scaleFactors[3729] = 0.0;
scaleFactors[3728] = 0.0;
scaleFactors[3727] = 0.0;
scaleFactors[3726] = 0.0;
scaleFactors[3725] = 0.0;
scaleFactors[3724] = 0.0;
scaleFactors[3723] = 0.0;
scaleFactors[3722] = 0.0;
scaleFactors[3721] = 0.0;
scaleFactors[3720] = 0.0;
scaleFactors[3719] = 0.0;
scaleFactors[3718] = 0.0;
scaleFactors[3717] = 0.0;
scaleFactors[3716] = 0.0;
scaleFactors[3715] = 0.0;
scaleFactors[3714] = 0.0;
scaleFactors[3713] = 0.0;
scaleFactors[3712] = 0.0;
scaleFactors[3711] = 0.0;
scaleFactors[3710] = 0.0;
scaleFactors[3709] = 0.0;
scaleFactors[3708] = 0.0;
scaleFactors[3707] = 0.0;
scaleFactors[3706] = 0.0;
scaleFactors[3705] = 0.0;
scaleFactors[3704] = 0.0;
scaleFactors[3703] = 0.0;
scaleFactors[3702] = 0.0;
scaleFactors[3701] = 0.0;
scaleFactors[3700] = 0.0;
scaleFactors[3699] = 0.0;
scaleFactors[3698] = 0.0;
scaleFactors[3697] = 0.0;
scaleFactors[3696] = 0.0;
scaleFactors[3695] = 0.0;
scaleFactors[3694] = 0.0;
scaleFactors[3693] = 0.0;
scaleFactors[3692] = 0.0;
scaleFactors[3691] = 0.0;
scaleFactors[3690] = 0.0;
scaleFactors[3689] = 0.0;
scaleFactors[3688] = 0.0;
scaleFactors[3687] = 0.0;
scaleFactors[3686] = 0.0;
scaleFactors[3685] = 0.0;
scaleFactors[3684] = 0.0;
scaleFactors[3683] = 0.0;
scaleFactors[3682] = 0.0;
scaleFactors[3681] = 0.0;
scaleFactors[3680] = 0.0;
scaleFactors[3679] = 0.0;
scaleFactors[3678] = 0.0;
scaleFactors[3677] = 0.0;
scaleFactors[3676] = 0.0;
scaleFactors[3675] = 0.0;
scaleFactors[3674] = 0.0;
scaleFactors[3673] = 0.0;
scaleFactors[3672] = 0.0;
scaleFactors[3671] = 0.0;
scaleFactors[3670] = 0.0;
scaleFactors[3669] = 0.0;
scaleFactors[3668] = 0.0;
scaleFactors[3667] = 0.0;
scaleFactors[3666] = 0.0;
scaleFactors[3665] = 0.0;
scaleFactors[3664] = 0.0;
scaleFactors[3663] = 0.0;
scaleFactors[3662] = 0.0;
scaleFactors[3661] = 0.0;
scaleFactors[3660] = 0.0;
scaleFactors[3659] = 0.0;
scaleFactors[3658] = 0.0;
scaleFactors[3657] = 0.0;
scaleFactors[3656] = 0.0;
scaleFactors[3655] = 0.0;
scaleFactors[3654] = 0.0;
scaleFactors[3653] = 0.0;
scaleFactors[3652] = 0.0;
scaleFactors[3651] = 0.0;
scaleFactors[3650] = 0.0;
scaleFactors[3649] = 0.0;
scaleFactors[3648] = 0.0;
scaleFactors[3647] = 0.0;
scaleFactors[3646] = 0.0;
scaleFactors[3645] = 0.0;
scaleFactors[3644] = 0.0;
scaleFactors[3643] = 0.0;
scaleFactors[3642] = 0.0;
scaleFactors[3641] = 0.0;
scaleFactors[3640] = 0.0;
scaleFactors[3639] = 0.0;
scaleFactors[3638] = 0.0;
scaleFactors[3637] = 0.0;
scaleFactors[3636] = 0.0;
scaleFactors[3635] = 0.0;
scaleFactors[3634] = 0.0;
scaleFactors[3633] = 0.0;
scaleFactors[3632] = 0.0;
scaleFactors[3631] = 0.0;
scaleFactors[3630] = 0.0;
scaleFactors[3629] = 0.0;
scaleFactors[3628] = 0.0;
scaleFactors[3627] = 0.0;
scaleFactors[3626] = 0.0;
scaleFactors[3625] = 0.0;
scaleFactors[3624] = 0.0;
scaleFactors[3623] = 0.0;
scaleFactors[3622] = 0.0;
scaleFactors[3621] = 0.0;
scaleFactors[3620] = 0.0;
scaleFactors[3619] = 0.0;
scaleFactors[3618] = 0.0;
scaleFactors[3617] = 0.0;
scaleFactors[3616] = 0.0;
scaleFactors[3615] = 0.0;
scaleFactors[3614] = 0.0;
scaleFactors[3613] = 0.0;
scaleFactors[3612] = 0.0;
scaleFactors[3611] = 0.0;
scaleFactors[3610] = 0.0;
scaleFactors[3609] = 0.0;
scaleFactors[3608] = 0.0;
scaleFactors[3607] = 0.0;
scaleFactors[3606] = 0.0;
scaleFactors[3605] = 0.0;
scaleFactors[3604] = 0.0;
scaleFactors[3603] = 0.0;
scaleFactors[3602] = 0.0;
scaleFactors[3601] = 0.0;
scaleFactors[3600] = 0.0;
scaleFactors[3599] = 0.0;
scaleFactors[3598] = 0.0;
scaleFactors[3597] = 0.0;
scaleFactors[3596] = 0.0;
scaleFactors[3595] = 0.0;
scaleFactors[3594] = 0.0;
scaleFactors[3593] = 0.0;
scaleFactors[3592] = 0.0;
scaleFactors[3591] = 0.0;
scaleFactors[3590] = 0.0;
scaleFactors[3589] = 0.0;
scaleFactors[3588] = 0.0;
scaleFactors[3587] = 0.0;
scaleFactors[3586] = 0.0;
scaleFactors[3585] = 0.0;
scaleFactors[3584] = 0.0;
scaleFactors[3583] = 0.0;
scaleFactors[3582] = 0.0;
scaleFactors[3581] = 0.0;
scaleFactors[3580] = 0.0;
scaleFactors[3579] = 0.0;
scaleFactors[3578] = 0.0;
scaleFactors[3577] = 0.0;
scaleFactors[3576] = 0.0;
scaleFactors[3575] = 0.0;
scaleFactors[3574] = 0.0;
scaleFactors[3573] = 0.0;
scaleFactors[3572] = 0.0;
scaleFactors[3571] = 0.0;
scaleFactors[3570] = 0.0;
scaleFactors[3569] = 0.0;
scaleFactors[3568] = 0.0;
scaleFactors[3567] = 0.0;
scaleFactors[3566] = 0.0;
scaleFactors[3565] = 0.0;
scaleFactors[3564] = 0.0;
scaleFactors[3563] = 0.0;
scaleFactors[3562] = 0.0;
scaleFactors[3561] = 0.0;
scaleFactors[3560] = 0.0;
scaleFactors[3559] = 0.0;
scaleFactors[3558] = 0.0;
scaleFactors[3557] = 0.0;
scaleFactors[3556] = 0.0;
scaleFactors[3555] = 0.0;
scaleFactors[3554] = 0.0;
scaleFactors[3553] = 0.0;
scaleFactors[3552] = 0.0;
scaleFactors[3551] = 0.0;
scaleFactors[3550] = 0.0;
scaleFactors[3549] = 0.0;
scaleFactors[3548] = 0.0;
scaleFactors[3547] = 0.0;
scaleFactors[3546] = 0.0;
scaleFactors[3545] = 0.0;
scaleFactors[3544] = 0.0;
scaleFactors[3543] = 0.0;
scaleFactors[3542] = 0.0;
scaleFactors[3541] = 0.0;
scaleFactors[3540] = 0.0;
scaleFactors[3539] = 0.0;
scaleFactors[3538] = 0.0;
scaleFactors[3537] = 0.0;
scaleFactors[3536] = 0.0;
scaleFactors[3535] = 0.0;
scaleFactors[3534] = 0.0;
scaleFactors[3533] = 0.0;
scaleFactors[3532] = 0.0;
scaleFactors[3531] = 0.0;
scaleFactors[3530] = 0.0;
scaleFactors[3529] = 0.0;
scaleFactors[3528] = 0.0;
scaleFactors[3527] = 0.0;
scaleFactors[3526] = 0.0;
scaleFactors[3525] = 0.0;
scaleFactors[3524] = 0.0;
scaleFactors[3523] = 0.0;
scaleFactors[3522] = 0.0;
scaleFactors[3521] = 0.0;
scaleFactors[3520] = 0.0;
scaleFactors[3519] = 0.0;
scaleFactors[3518] = 0.0;
scaleFactors[3517] = 0.0;
scaleFactors[3516] = 0.0;
scaleFactors[3515] = 0.0;
scaleFactors[3514] = 0.0;
scaleFactors[3513] = 0.0;
scaleFactors[3512] = 0.0;
scaleFactors[3511] = 0.0;
scaleFactors[3510] = 0.0;
scaleFactors[3509] = 0.0;
scaleFactors[3508] = 0.0;
scaleFactors[3507] = 0.0;
scaleFactors[3506] = 0.0;
scaleFactors[3505] = 0.0;
scaleFactors[3504] = 0.0;
scaleFactors[3503] = 0.0;
scaleFactors[3502] = 0.0;
scaleFactors[3501] = 0.0;
scaleFactors[3500] = 0.0;
scaleFactors[3499] = 0.0;
scaleFactors[3498] = 0.0;
scaleFactors[3497] = 0.0;
scaleFactors[3496] = 0.0;
scaleFactors[3495] = 0.0;
scaleFactors[3494] = 0.0;
scaleFactors[3493] = 0.0;
scaleFactors[3492] = 0.0;
scaleFactors[3491] = 0.0;
scaleFactors[3490] = 0.0;
scaleFactors[3489] = 0.0;
scaleFactors[3488] = 0.0;
scaleFactors[3487] = 0.0;
scaleFactors[3486] = 0.0;
scaleFactors[3485] = 0.0;
scaleFactors[3484] = 0.0;
scaleFactors[3483] = 0.0;
scaleFactors[3482] = 0.0;
scaleFactors[3481] = 0.0;
scaleFactors[3480] = 0.0;
scaleFactors[3479] = 0.0;
scaleFactors[3478] = 0.0;
scaleFactors[3477] = 0.0;
scaleFactors[3476] = 0.0;
scaleFactors[3475] = 0.0;
scaleFactors[3474] = 0.0;
scaleFactors[3473] = 0.0;
scaleFactors[3472] = 0.0;
scaleFactors[3471] = 0.0;
scaleFactors[3470] = 0.0;
scaleFactors[3469] = 0.0;
scaleFactors[3468] = 0.0;
scaleFactors[3467] = 0.0;
scaleFactors[3466] = 0.0;
scaleFactors[3465] = 0.0;
scaleFactors[3464] = 0.0;
scaleFactors[3463] = 0.0;
scaleFactors[3462] = 0.0;
scaleFactors[3461] = 0.0;
scaleFactors[3460] = 0.0;
scaleFactors[3459] = 0.0;
scaleFactors[3458] = 0.0;
scaleFactors[3457] = 0.0;
scaleFactors[3456] = 0.0;
scaleFactors[3455] = 0.0;
scaleFactors[3454] = 0.0;
scaleFactors[3453] = 0.0;
scaleFactors[3452] = 0.0;
scaleFactors[3451] = 0.0;
scaleFactors[3450] = 0.0;
scaleFactors[3449] = 0.0;
scaleFactors[3448] = 0.0;
scaleFactors[3447] = 0.0;
scaleFactors[3446] = 0.0;
scaleFactors[3445] = 0.0;
scaleFactors[3444] = 0.0;
scaleFactors[3443] = 0.0;
scaleFactors[3442] = 0.0;
scaleFactors[3441] = 0.0;
scaleFactors[3440] = 0.0;
scaleFactors[3439] = 0.0;
scaleFactors[3438] = 0.0;
scaleFactors[3437] = 0.0;
scaleFactors[3436] = 0.0;
scaleFactors[3435] = 0.0;
scaleFactors[3434] = 0.0;
scaleFactors[3433] = 0.0;
scaleFactors[3432] = 0.0;
scaleFactors[3431] = 0.0;
scaleFactors[3430] = 0.0;
scaleFactors[3429] = 0.0;
scaleFactors[3428] = 0.0;
scaleFactors[3427] = 0.0;
scaleFactors[3426] = 0.0;
scaleFactors[3425] = 0.0;
scaleFactors[3424] = 0.0;
scaleFactors[3423] = 0.0;
scaleFactors[3422] = 0.0;
scaleFactors[3421] = 0.0;
scaleFactors[3420] = 0.0;
scaleFactors[3419] = 0.0;
scaleFactors[3418] = 0.0;
scaleFactors[3417] = 0.0;
scaleFactors[3416] = 0.0;
scaleFactors[3415] = 0.0;
scaleFactors[3414] = 0.0;
scaleFactors[3413] = 0.0;
scaleFactors[3412] = 0.0;
scaleFactors[3411] = 0.0;
scaleFactors[3410] = 0.0;
scaleFactors[3409] = 0.0;
scaleFactors[3408] = 0.0;
scaleFactors[3407] = 0.0;
scaleFactors[3406] = 0.0;
scaleFactors[3405] = 0.0;
scaleFactors[3404] = 0.0;
scaleFactors[3403] = 0.0;
scaleFactors[3402] = 0.0;
scaleFactors[3401] = 0.0;
scaleFactors[3400] = 0.0;
scaleFactors[3399] = 0.0;
scaleFactors[3398] = 0.0;
scaleFactors[3397] = 0.0;
scaleFactors[3396] = 0.0;
scaleFactors[3395] = 0.0;
scaleFactors[3394] = 0.0;
scaleFactors[3393] = 0.0;
scaleFactors[3392] = 0.0;
scaleFactors[3391] = 0.0;
scaleFactors[3390] = 0.0;
scaleFactors[3389] = 0.0;
scaleFactors[3388] = 0.0;
scaleFactors[3387] = 0.0;
scaleFactors[3386] = 0.0;
scaleFactors[3385] = 0.0;
scaleFactors[3384] = 0.0;
scaleFactors[3383] = 0.0;
scaleFactors[3382] = 0.0;
scaleFactors[3381] = 0.0;
scaleFactors[3380] = 0.0;
scaleFactors[3379] = 0.0;
scaleFactors[3378] = 0.0;
scaleFactors[3377] = 0.0;
scaleFactors[3376] = 0.0;
scaleFactors[3375] = 0.0;
scaleFactors[3374] = 0.0;
scaleFactors[3373] = 0.0;
scaleFactors[3372] = 0.0;
scaleFactors[3371] = 0.0;
scaleFactors[3370] = 0.0;
scaleFactors[3369] = 0.0;
scaleFactors[3368] = 0.0;
scaleFactors[3367] = 0.0;
scaleFactors[3366] = 0.0;
scaleFactors[3365] = 0.0;
scaleFactors[3364] = 0.0;
scaleFactors[3363] = 0.0;
scaleFactors[3362] = 0.0;
scaleFactors[3361] = 0.0;
scaleFactors[3360] = 0.0;
scaleFactors[3359] = 0.0;
scaleFactors[3358] = 0.0;
scaleFactors[3357] = 0.0;
scaleFactors[3356] = 0.0;
scaleFactors[3355] = 0.0;
scaleFactors[3354] = 0.0;
scaleFactors[3353] = 0.0;
scaleFactors[3352] = 0.0;
scaleFactors[3351] = 0.0;
scaleFactors[3350] = 0.0;
scaleFactors[3349] = 0.0;
scaleFactors[3348] = 0.0;
scaleFactors[3347] = 0.0;
scaleFactors[3346] = 0.0;
scaleFactors[3345] = 0.0;
scaleFactors[3344] = 0.0;
scaleFactors[3343] = 0.0;
scaleFactors[3342] = 0.0;
scaleFactors[3341] = 0.0;
scaleFactors[3340] = 0.0;
scaleFactors[3339] = 0.0;
scaleFactors[3338] = 0.0;
scaleFactors[3337] = 0.0;
scaleFactors[3336] = 0.0;
scaleFactors[3335] = 0.0;
scaleFactors[3334] = 0.0;
scaleFactors[3333] = 0.0;
scaleFactors[3332] = 0.0;
scaleFactors[3331] = 0.0;
scaleFactors[3330] = 0.0;
scaleFactors[3329] = 0.0;
scaleFactors[3328] = 0.0;
scaleFactors[3327] = 0.0;
scaleFactors[3326] = 0.0;
scaleFactors[3325] = 0.0;
scaleFactors[3324] = 0.0;
scaleFactors[3323] = 0.0;
scaleFactors[3322] = 0.0;
scaleFactors[3321] = 0.0;
scaleFactors[3320] = 0.0;
scaleFactors[3319] = 0.0;
scaleFactors[3318] = 0.0;
scaleFactors[3317] = 0.0;
scaleFactors[3316] = 0.0;
scaleFactors[3315] = 0.0;
scaleFactors[3314] = 0.0;
scaleFactors[3313] = 0.0;
scaleFactors[3312] = 0.0;
scaleFactors[3311] = 0.0;
scaleFactors[3310] = 0.0;
scaleFactors[3309] = 0.0;
scaleFactors[3308] = 0.0;
scaleFactors[3307] = 0.0;
scaleFactors[3306] = 0.0;
scaleFactors[3305] = 0.0;
scaleFactors[3304] = 0.0;
scaleFactors[3303] = 0.0;
scaleFactors[3302] = 0.0;
scaleFactors[3301] = 0.0;
scaleFactors[3300] = 0.0;
scaleFactors[3299] = 0.0;
scaleFactors[3298] = 0.0;
scaleFactors[3297] = 0.0;
scaleFactors[3296] = 0.0;
scaleFactors[3295] = 0.0;
scaleFactors[3294] = 0.0;
scaleFactors[3293] = 0.0;
scaleFactors[3292] = 0.0;
scaleFactors[3291] = 0.0;
scaleFactors[3290] = 0.0;
scaleFactors[3289] = 0.0;
scaleFactors[3288] = 0.0;
scaleFactors[3287] = 0.0;
scaleFactors[3286] = 0.0;
scaleFactors[3285] = 0.0;
scaleFactors[3284] = 0.0;
scaleFactors[3283] = 0.0;
scaleFactors[3282] = 0.0;
scaleFactors[3281] = 0.0;
scaleFactors[3280] = 0.0;
scaleFactors[3279] = 0.0;
scaleFactors[3278] = 0.0;
scaleFactors[3277] = 0.0;
scaleFactors[3276] = 0.0;
scaleFactors[3275] = 0.0;
scaleFactors[3274] = 0.0;
scaleFactors[3273] = 0.0;
scaleFactors[3272] = 0.0;
scaleFactors[3271] = 0.0;
scaleFactors[3270] = 0.0;
scaleFactors[3269] = 0.0;
scaleFactors[3268] = 0.0;
scaleFactors[3267] = 0.0;
scaleFactors[3266] = 0.0;
scaleFactors[3265] = 0.0;
scaleFactors[3264] = 0.0;
scaleFactors[3263] = 0.0;
scaleFactors[3262] = 0.0;
scaleFactors[3261] = 0.0;
scaleFactors[3260] = 0.0;
scaleFactors[3259] = 0.0;
scaleFactors[3258] = 0.0;
scaleFactors[3257] = 0.0;
scaleFactors[3256] = 0.0;
scaleFactors[3255] = 0.0;
scaleFactors[3254] = 0.0;
scaleFactors[3253] = 0.0;
scaleFactors[3252] = 0.0;
scaleFactors[3251] = 0.0;
scaleFactors[3250] = 0.0;
scaleFactors[3249] = 0.0;
scaleFactors[3248] = 0.0;
scaleFactors[3247] = 0.0;
scaleFactors[3246] = 0.0;
scaleFactors[3245] = 0.0;
scaleFactors[3244] = 0.0;
scaleFactors[3243] = 0.0;
scaleFactors[3242] = 0.0;
scaleFactors[3241] = 0.0;
scaleFactors[3240] = 0.0;
scaleFactors[3239] = 0.0;
scaleFactors[3238] = 0.0;
scaleFactors[3237] = 0.0;
scaleFactors[3236] = 0.0;
scaleFactors[3235] = 0.0;
scaleFactors[3234] = 0.0;
scaleFactors[3233] = 0.0;
scaleFactors[3232] = 0.0;
scaleFactors[3231] = 0.0;
scaleFactors[3230] = 0.0;
scaleFactors[3229] = 0.0;
scaleFactors[3228] = 0.0;
scaleFactors[3227] = 0.0;
scaleFactors[3226] = 0.0;
scaleFactors[3225] = 0.0;
scaleFactors[3224] = 0.0;
scaleFactors[3223] = 0.0;
scaleFactors[3222] = 0.0;
scaleFactors[3221] = 0.0;
scaleFactors[3220] = 0.0;
scaleFactors[3219] = 0.0;
scaleFactors[3218] = 0.0;
scaleFactors[3217] = 0.0;
scaleFactors[3216] = 0.0;
scaleFactors[3215] = 0.0;
scaleFactors[3214] = 0.0;
scaleFactors[3213] = 0.0;
scaleFactors[3212] = 0.0;
scaleFactors[3211] = 0.0;
scaleFactors[3210] = 0.0;
scaleFactors[3209] = 0.0;
scaleFactors[3208] = 0.0;
scaleFactors[3207] = 0.0;
scaleFactors[3206] = 0.0;
scaleFactors[3205] = 0.0;
scaleFactors[3204] = 0.0;
scaleFactors[3203] = 0.0;
scaleFactors[3202] = 0.0;
scaleFactors[3201] = 0.0;
scaleFactors[3200] = 0.0;
scaleFactors[3199] = 0.0;
scaleFactors[3198] = 0.0;
scaleFactors[3197] = 0.0;
scaleFactors[3196] = 0.0;
scaleFactors[3195] = 0.0;
scaleFactors[3194] = 0.0;
scaleFactors[3193] = 0.0;
scaleFactors[3192] = 0.0;
scaleFactors[3191] = 0.0;
scaleFactors[3190] = 0.0;
scaleFactors[3189] = 0.0;
scaleFactors[3188] = 0.0;
scaleFactors[3187] = 0.0;
scaleFactors[3186] = 0.0;
scaleFactors[3185] = 0.0;
scaleFactors[3184] = 0.0;
scaleFactors[3183] = 0.0;
scaleFactors[3182] = 0.0;
scaleFactors[3181] = 0.0;
scaleFactors[3180] = 0.0;
scaleFactors[3179] = 0.0;
scaleFactors[3178] = 0.0;
scaleFactors[3177] = 0.0;
scaleFactors[3176] = 0.0;
scaleFactors[3175] = 0.0;
scaleFactors[3174] = 0.0;
scaleFactors[3173] = 0.0;
scaleFactors[3172] = 0.0;
scaleFactors[3171] = 0.0;
scaleFactors[3170] = 0.0;
scaleFactors[3169] = 0.0;
scaleFactors[3168] = 0.0;
scaleFactors[3167] = 0.0;
scaleFactors[3166] = 0.0;
scaleFactors[3165] = 0.0;
scaleFactors[3164] = 0.0;
scaleFactors[3163] = 0.0;
scaleFactors[3162] = 0.0;
scaleFactors[3161] = 0.0;
scaleFactors[3160] = 0.0;
scaleFactors[3159] = 0.0;
scaleFactors[3158] = 0.0;
scaleFactors[3157] = 0.0;
scaleFactors[3156] = 0.0;
scaleFactors[3155] = 0.0;
scaleFactors[3154] = 0.0;
scaleFactors[3153] = 0.0;
scaleFactors[3152] = 0.0;
scaleFactors[3151] = 0.0;
scaleFactors[3150] = 0.0;
scaleFactors[3149] = 0.0;
scaleFactors[3148] = 0.0;
scaleFactors[3147] = 0.0;
scaleFactors[3146] = 0.0;
scaleFactors[3145] = 0.0;
scaleFactors[3144] = 0.0;
scaleFactors[3143] = 0.0;
scaleFactors[3142] = 0.0;
scaleFactors[3141] = 0.0;
scaleFactors[3140] = 0.0;
scaleFactors[3139] = 0.0;
scaleFactors[3138] = 0.0;
scaleFactors[3137] = 0.0;
scaleFactors[3136] = 0.0;
scaleFactors[3135] = 0.0;
scaleFactors[3134] = 0.0;
scaleFactors[3133] = 0.0;
scaleFactors[3132] = 0.0;
scaleFactors[3131] = 0.0;
scaleFactors[3130] = 0.0;
scaleFactors[3129] = 0.0;
scaleFactors[3128] = 0.0;
scaleFactors[3127] = 0.0;
scaleFactors[3126] = 0.0;
scaleFactors[3125] = 0.0;
scaleFactors[3124] = 0.0;
scaleFactors[3123] = 0.0;
scaleFactors[3122] = 0.0;
scaleFactors[3121] = 0.0;
scaleFactors[3120] = 0.0;
scaleFactors[3119] = 0.0;
scaleFactors[3118] = 0.0;
scaleFactors[3117] = 0.0;
scaleFactors[3116] = 0.0;
scaleFactors[3115] = 0.0;
scaleFactors[3114] = 0.0;
scaleFactors[3113] = 0.0;
scaleFactors[3112] = 0.0;
scaleFactors[3111] = 0.0;
scaleFactors[3110] = 0.0;
scaleFactors[3109] = 0.0;
scaleFactors[3108] = 0.0;
scaleFactors[3107] = 0.0;
scaleFactors[3106] = 0.0;
scaleFactors[3105] = 0.0;
scaleFactors[3104] = 0.0;
scaleFactors[3103] = 0.0;
scaleFactors[3102] = 0.0;
scaleFactors[3101] = 0.0;
scaleFactors[3100] = 0.0;
scaleFactors[3099] = 0.0;
scaleFactors[3098] = 0.0;
scaleFactors[3097] = 0.0;
scaleFactors[3096] = 0.0;
scaleFactors[3095] = 0.0;
scaleFactors[3094] = 0.0;
scaleFactors[3093] = 0.0;
scaleFactors[3092] = 0.0;
scaleFactors[3091] = 0.0;
scaleFactors[3090] = 0.0;
scaleFactors[3089] = 0.0;
scaleFactors[3088] = 0.0;
scaleFactors[3087] = 0.0;
scaleFactors[3086] = 0.0;
scaleFactors[3085] = 0.0;
scaleFactors[3084] = 0.0;
scaleFactors[3083] = 0.0;
scaleFactors[3082] = 0.0;
scaleFactors[3081] = 0.0;
scaleFactors[3080] = 0.0;
scaleFactors[3079] = 0.0;
scaleFactors[3078] = 0.0;
scaleFactors[3077] = 0.0;
scaleFactors[3076] = 0.0;
scaleFactors[3075] = 0.0;
scaleFactors[3074] = 0.0;
scaleFactors[3073] = 0.0;
scaleFactors[3072] = 0.0;
scaleFactors[3071] = 0.0;
scaleFactors[3070] = 0.0;
scaleFactors[3069] = 0.0;
scaleFactors[3068] = 0.0;
scaleFactors[3067] = 0.0;
scaleFactors[3066] = 0.0;
scaleFactors[3065] = 0.0;
scaleFactors[3064] = 0.0;
scaleFactors[3063] = 0.0;
scaleFactors[3062] = 0.0;
scaleFactors[3061] = 0.0;
scaleFactors[3060] = 0.0;
scaleFactors[3059] = 0.0;
scaleFactors[3058] = 0.0;
scaleFactors[3057] = 0.0;
scaleFactors[3056] = 0.0;
scaleFactors[3055] = 0.0;
scaleFactors[3054] = 0.0;
scaleFactors[3053] = 0.0;
scaleFactors[3052] = 0.0;
scaleFactors[3051] = 0.0;
scaleFactors[3050] = 0.0;
scaleFactors[3049] = 0.0;
scaleFactors[3048] = 0.0;
scaleFactors[3047] = 0.0;
scaleFactors[3046] = 0.0;
scaleFactors[3045] = 0.0;
scaleFactors[3044] = 0.0;
scaleFactors[3043] = 0.0;
scaleFactors[3042] = 0.0;
scaleFactors[3041] = 0.0;
scaleFactors[3040] = 0.0;
scaleFactors[3039] = 0.0;
scaleFactors[3038] = 0.0;
scaleFactors[3037] = 0.0;
scaleFactors[3036] = 0.0;
scaleFactors[3035] = 0.0;
scaleFactors[3034] = 0.0;
scaleFactors[3033] = 0.0;
scaleFactors[3032] = 0.0;
scaleFactors[3031] = 0.0;
scaleFactors[3030] = 0.0;
scaleFactors[3029] = 0.0;
scaleFactors[3028] = 0.0;
scaleFactors[3027] = 0.0;
scaleFactors[3026] = 0.0;
scaleFactors[3025] = 0.0;
scaleFactors[3024] = 0.0;
scaleFactors[3023] = 0.0;
scaleFactors[3022] = 0.0;
scaleFactors[3021] = 0.0;
scaleFactors[3020] = 0.0;
scaleFactors[3019] = 0.0;
scaleFactors[3018] = 0.0;
scaleFactors[3017] = 0.0;
scaleFactors[3016] = 0.0;
scaleFactors[3015] = 0.0;
scaleFactors[3014] = 0.0;
scaleFactors[3013] = 0.0;
scaleFactors[3012] = 0.0;
scaleFactors[3011] = 0.0;
scaleFactors[3010] = 0.0;
scaleFactors[3009] = 0.0;
scaleFactors[3008] = 0.0;
scaleFactors[3007] = 0.0;
scaleFactors[3006] = 0.0;
scaleFactors[3005] = 0.0;
scaleFactors[3004] = 0.0;
scaleFactors[3003] = 0.0;
scaleFactors[3002] = 0.0;
scaleFactors[3001] = 0.0;
scaleFactors[3000] = 0.0;
scaleFactors[2999] = 0.0;
scaleFactors[2998] = 0.0;
scaleFactors[2997] = 0.0;
scaleFactors[2996] = 0.0;
scaleFactors[2995] = 0.0;
scaleFactors[2994] = 0.0;
scaleFactors[2993] = 0.0;
scaleFactors[2992] = 0.0;
scaleFactors[2991] = 0.0;
scaleFactors[2990] = 0.0;
scaleFactors[2989] = 0.0;
scaleFactors[2988] = 0.0;
scaleFactors[2987] = 0.0;
scaleFactors[2986] = 0.0;
scaleFactors[2985] = 0.0;
scaleFactors[2984] = 0.0;
scaleFactors[2983] = 0.0;
scaleFactors[2982] = 0.0;
scaleFactors[2981] = 0.0;
scaleFactors[2980] = 0.0;
scaleFactors[2979] = 0.0;
scaleFactors[2978] = 0.0;
scaleFactors[2977] = 0.0;
scaleFactors[2976] = 0.0;
scaleFactors[2975] = 0.0;
scaleFactors[2974] = 0.0;
scaleFactors[2973] = 0.0;
scaleFactors[2972] = 0.0;
scaleFactors[2971] = 0.0;
scaleFactors[2970] = 0.0;
scaleFactors[2969] = 0.0;
scaleFactors[2968] = 0.0;
scaleFactors[2967] = 0.0;
scaleFactors[2966] = 0.0;
scaleFactors[2965] = 0.0;
scaleFactors[2964] = 0.0;
scaleFactors[2963] = 0.0;
scaleFactors[2962] = 0.0;
scaleFactors[2961] = 0.0;
scaleFactors[2960] = 0.0;
scaleFactors[2959] = 0.0;
scaleFactors[2958] = 0.0;
scaleFactors[2957] = 0.0;
scaleFactors[2956] = 0.0;
scaleFactors[2955] = 0.0;
scaleFactors[2954] = 0.0;
scaleFactors[2953] = 0.0;
scaleFactors[2952] = 0.0;
scaleFactors[2951] = 0.0;
scaleFactors[2950] = 0.0;
scaleFactors[2949] = 0.0;
scaleFactors[2948] = 0.0;
scaleFactors[2947] = 0.0;
scaleFactors[2946] = 0.0;
scaleFactors[2945] = 0.0;
scaleFactors[2944] = 0.0;
scaleFactors[2943] = 0.0;
scaleFactors[2942] = 0.0;
scaleFactors[2941] = 0.0;
scaleFactors[2940] = 0.0;
scaleFactors[2939] = 0.0;
scaleFactors[2938] = 0.0;
scaleFactors[2937] = 0.0;
scaleFactors[2936] = 0.0;
scaleFactors[2935] = 0.0;
scaleFactors[2934] = 0.0;
scaleFactors[2933] = 0.0;
scaleFactors[2932] = 0.0;
scaleFactors[2931] = 0.0;
scaleFactors[2930] = 0.0;
scaleFactors[2929] = 0.0;
scaleFactors[2928] = 0.0;
scaleFactors[2927] = 0.0;
scaleFactors[2926] = 0.0;
scaleFactors[2925] = 0.0;
scaleFactors[2924] = 0.0;
scaleFactors[2923] = 0.0;
scaleFactors[2922] = 0.0;
scaleFactors[2921] = 0.0;
scaleFactors[2920] = 0.0;
scaleFactors[2919] = 0.0;
scaleFactors[2918] = 0.0;
scaleFactors[2917] = 0.0;
scaleFactors[2916] = 0.0;
scaleFactors[2915] = 0.0;
scaleFactors[2914] = 0.0;
scaleFactors[2913] = 0.0;
scaleFactors[2912] = 0.0;
scaleFactors[2911] = 0.0;
scaleFactors[2910] = 0.0;
scaleFactors[2909] = 0.0;
scaleFactors[2908] = 0.0;
scaleFactors[2907] = 0.0;
scaleFactors[2906] = 0.0;
scaleFactors[2905] = 0.0;
scaleFactors[2904] = 0.0;
scaleFactors[2903] = 0.0;
scaleFactors[2902] = 0.0;
scaleFactors[2901] = 0.0;
scaleFactors[2900] = 0.0;
scaleFactors[2899] = 0.0;
scaleFactors[2898] = 0.0;
scaleFactors[2897] = 0.0;
scaleFactors[2896] = 0.0;
scaleFactors[2895] = 0.0;
scaleFactors[2894] = 0.0;
scaleFactors[2893] = 0.0;
scaleFactors[2892] = 0.0;
scaleFactors[2891] = 0.0;
scaleFactors[2890] = 0.0;
scaleFactors[2889] = 0.0;
scaleFactors[2888] = 0.0;
scaleFactors[2887] = 0.0;
scaleFactors[2886] = 0.0;
scaleFactors[2885] = 0.0;
scaleFactors[2884] = 0.0;
scaleFactors[2883] = 0.0;
scaleFactors[2882] = 0.0;
scaleFactors[2881] = 0.0;
scaleFactors[2880] = 0.0;
scaleFactors[2879] = 0.0;
scaleFactors[2878] = 0.0;
scaleFactors[2877] = 0.0;
scaleFactors[2876] = 0.0;
scaleFactors[2875] = 0.0;
scaleFactors[2874] = 0.0;
scaleFactors[2873] = 0.0;
scaleFactors[2872] = 0.0;
scaleFactors[2871] = 0.0;
scaleFactors[2870] = 0.0;
scaleFactors[2869] = 0.0;
scaleFactors[2868] = 0.0;
scaleFactors[2867] = 0.0;
scaleFactors[2866] = 0.0;
scaleFactors[2865] = 0.0;
scaleFactors[2864] = 0.0;
scaleFactors[2863] = 0.0;
scaleFactors[2862] = 0.0;
scaleFactors[2861] = 0.0;
scaleFactors[2860] = 0.0;
scaleFactors[2859] = 0.0;
scaleFactors[2858] = 0.0;
scaleFactors[2857] = 0.0;
scaleFactors[2856] = 0.0;
scaleFactors[2855] = 0.0;
scaleFactors[2854] = 0.0;
scaleFactors[2853] = 0.0;
scaleFactors[2852] = 0.0;
scaleFactors[2851] = 0.0;
scaleFactors[2850] = 0.0;
scaleFactors[2849] = 0.0;
scaleFactors[2848] = 0.0;
scaleFactors[2847] = 0.0;
scaleFactors[2846] = 0.0;
scaleFactors[2845] = 0.0;
scaleFactors[2844] = 0.0;
scaleFactors[2843] = 0.0;
scaleFactors[2842] = 0.0;
scaleFactors[2841] = 0.0;
scaleFactors[2840] = 0.0;
scaleFactors[2839] = 0.0;
scaleFactors[2838] = 0.0;
scaleFactors[2837] = 0.0;
scaleFactors[2836] = 0.0;
scaleFactors[2835] = 0.0;
scaleFactors[2834] = 0.0;
scaleFactors[2833] = 0.0;
scaleFactors[2832] = 0.0;
scaleFactors[2831] = 0.0;
scaleFactors[2830] = 0.0;
scaleFactors[2829] = 0.0;
scaleFactors[2828] = 0.0;
scaleFactors[2827] = 0.0;
scaleFactors[2826] = 0.0;
scaleFactors[2825] = 0.0;
scaleFactors[2824] = 0.0;
scaleFactors[2823] = 0.0;
scaleFactors[2822] = 0.0;
scaleFactors[2821] = 0.0;
scaleFactors[2820] = 0.0;
scaleFactors[2819] = 0.0;
scaleFactors[2818] = 0.0;
scaleFactors[2817] = 0.0;
scaleFactors[2816] = 0.0;
scaleFactors[2815] = 0.0;
scaleFactors[2814] = 0.0;
scaleFactors[2813] = 0.0;
scaleFactors[2812] = 0.0;
scaleFactors[2811] = 0.0;
scaleFactors[2810] = 0.0;
scaleFactors[2809] = 0.0;
scaleFactors[2808] = 0.0;
scaleFactors[2807] = 0.0;
scaleFactors[2806] = 0.0;
scaleFactors[2805] = 0.0;
scaleFactors[2804] = 0.0;
scaleFactors[2803] = 0.0;
scaleFactors[2802] = 0.0;
scaleFactors[2801] = 0.0;
scaleFactors[2800] = 0.0;
scaleFactors[2799] = 0.0;
scaleFactors[2798] = 0.0;
scaleFactors[2797] = 0.0;
scaleFactors[2796] = 0.0;
scaleFactors[2795] = 0.0;
scaleFactors[2794] = 0.0;
scaleFactors[2793] = 0.0;
scaleFactors[2792] = 0.0;
scaleFactors[2791] = 0.0;
scaleFactors[2790] = 0.0;
scaleFactors[2789] = 0.0;
scaleFactors[2788] = 0.0;
scaleFactors[2787] = 0.0;
scaleFactors[2786] = 0.0;
scaleFactors[2785] = 0.0;
scaleFactors[2784] = 0.0;
scaleFactors[2783] = 0.0;
scaleFactors[2782] = 0.0;
scaleFactors[2781] = 0.0;
scaleFactors[2780] = 0.0;
scaleFactors[2779] = 0.0;
scaleFactors[2778] = 0.0;
scaleFactors[2777] = 0.0;
scaleFactors[2776] = 0.0;
scaleFactors[2775] = 0.0;
scaleFactors[2774] = 0.0;
scaleFactors[2773] = 0.0;
scaleFactors[2772] = 0.0;
scaleFactors[2771] = 0.0;
scaleFactors[2770] = 0.0;
scaleFactors[2769] = 0.0;
scaleFactors[2768] = 0.0;
scaleFactors[2767] = 0.0;
scaleFactors[2766] = 0.0;
scaleFactors[2765] = 0.0;
scaleFactors[2764] = 0.0;
scaleFactors[2763] = 0.0;
scaleFactors[2762] = 0.0;
scaleFactors[2761] = 0.0;
scaleFactors[2760] = 0.0;
scaleFactors[2759] = 0.0;
scaleFactors[2758] = 0.0;
scaleFactors[2757] = 0.0;
scaleFactors[2756] = 0.0;
scaleFactors[2755] = 0.0;
scaleFactors[2754] = 0.0;
scaleFactors[2753] = 0.0;
scaleFactors[2752] = 0.0;
scaleFactors[2751] = 0.0;
scaleFactors[2750] = 0.0;
scaleFactors[2749] = 0.0;
scaleFactors[2748] = 0.0;
scaleFactors[2747] = 0.0;
scaleFactors[2746] = 0.0;
scaleFactors[2745] = 0.0;
scaleFactors[2744] = 0.0;
scaleFactors[2743] = 0.0;
scaleFactors[2742] = 0.0;
scaleFactors[2741] = 0.0;
scaleFactors[2740] = 0.0;
scaleFactors[2739] = 0.0;
scaleFactors[2738] = 0.0;
scaleFactors[2737] = 0.0;
scaleFactors[2736] = 0.0;
scaleFactors[2735] = 0.0;
scaleFactors[2734] = 0.0;
scaleFactors[2733] = 0.0;
scaleFactors[2732] = 0.0;
scaleFactors[2731] = 0.0;
scaleFactors[2730] = 0.0;
scaleFactors[2729] = 0.0;
scaleFactors[2728] = 0.0;
scaleFactors[2727] = 0.0;
scaleFactors[2726] = 0.0;
scaleFactors[2725] = 0.0;
scaleFactors[2724] = 0.0;
scaleFactors[2723] = 0.0;
scaleFactors[2722] = 0.0;
scaleFactors[2721] = 0.0;
scaleFactors[2720] = 0.0;
scaleFactors[2719] = 0.0;
scaleFactors[2718] = 0.0;
scaleFactors[2717] = 0.0;
scaleFactors[2716] = 0.0;
scaleFactors[2715] = 0.0;
scaleFactors[2714] = 0.0;
scaleFactors[2713] = 0.0;
scaleFactors[2712] = 0.0;
scaleFactors[2711] = 0.0;
scaleFactors[2710] = 0.0;
scaleFactors[2709] = 0.0;
scaleFactors[2708] = 0.0;
scaleFactors[2707] = 0.0;
scaleFactors[2706] = 0.0;
scaleFactors[2705] = 0.0;
scaleFactors[2704] = 0.0;
scaleFactors[2703] = 0.0;
scaleFactors[2702] = 0.0;
scaleFactors[2701] = 0.0;
scaleFactors[2700] = 0.0;
scaleFactors[2699] = 0.0;
scaleFactors[2698] = 0.0;
scaleFactors[2697] = 0.0;
scaleFactors[2696] = 0.0;
scaleFactors[2695] = 0.0;
scaleFactors[2694] = 0.0;
scaleFactors[2693] = 0.0;
scaleFactors[2692] = 0.0;
scaleFactors[2691] = 0.0;
scaleFactors[2690] = 0.0;
scaleFactors[2689] = 0.0;
scaleFactors[2688] = 0.0;
scaleFactors[2687] = 0.0;
scaleFactors[2686] = 0.0;
scaleFactors[2685] = 0.0;
scaleFactors[2684] = 0.0;
scaleFactors[2683] = 0.0;
scaleFactors[2682] = 0.0;
scaleFactors[2681] = 0.0;
scaleFactors[2680] = 0.0;
scaleFactors[2679] = 0.0;
scaleFactors[2678] = 0.0;
scaleFactors[2677] = 0.0;
scaleFactors[2676] = 0.0;
scaleFactors[2675] = 0.0;
scaleFactors[2674] = 0.0;
scaleFactors[2673] = 0.0;
scaleFactors[2672] = 0.0;
scaleFactors[2671] = 0.0;
scaleFactors[2670] = 0.0;
scaleFactors[2669] = 0.0;
scaleFactors[2668] = 0.0;
scaleFactors[2667] = 0.0;
scaleFactors[2666] = 0.0;
scaleFactors[2665] = 0.0;
scaleFactors[2664] = 0.0;
scaleFactors[2663] = 0.0;
scaleFactors[2662] = 0.0;
scaleFactors[2661] = 0.0;
scaleFactors[2660] = 0.0;
scaleFactors[2659] = 0.0;
scaleFactors[2658] = 0.0;
scaleFactors[2657] = 0.0;
scaleFactors[2656] = 0.0;
scaleFactors[2655] = 0.0;
scaleFactors[2654] = 0.0;
scaleFactors[2653] = 0.0;
scaleFactors[2652] = 0.0;
scaleFactors[2651] = 0.0;
scaleFactors[2650] = 0.0;
scaleFactors[2649] = 0.0;
scaleFactors[2648] = 0.0;
scaleFactors[2647] = 0.0;
scaleFactors[2646] = 0.0;
scaleFactors[2645] = 0.0;
scaleFactors[2644] = 0.0;
scaleFactors[2643] = 0.0;
scaleFactors[2642] = 0.0;
scaleFactors[2641] = 0.0;
scaleFactors[2640] = 0.0;
scaleFactors[2639] = 0.0;
scaleFactors[2638] = 0.0;
scaleFactors[2637] = 0.0;
scaleFactors[2636] = 0.0;
scaleFactors[2635] = 0.0;
scaleFactors[2634] = 0.0;
scaleFactors[2633] = 0.0;
scaleFactors[2632] = 0.0;
scaleFactors[2631] = 0.0;
scaleFactors[2630] = 0.0;
scaleFactors[2629] = 0.0;
scaleFactors[2628] = 0.0;
scaleFactors[2627] = 0.0;
scaleFactors[2626] = 0.0;
scaleFactors[2625] = 0.0;
scaleFactors[2624] = 0.0;
scaleFactors[2623] = 0.0;
scaleFactors[2622] = 0.0;
scaleFactors[2621] = 0.0;
scaleFactors[2620] = 0.0;
scaleFactors[2619] = 0.0;
scaleFactors[2618] = 0.0;
scaleFactors[2617] = 0.0;
scaleFactors[2616] = 0.0;
scaleFactors[2615] = 0.0;
scaleFactors[2614] = 0.0;
scaleFactors[2613] = 0.0;
scaleFactors[2612] = 0.0;
scaleFactors[2611] = 0.0;
scaleFactors[2610] = 0.0;
scaleFactors[2609] = 0.0;
scaleFactors[2608] = 0.0;
scaleFactors[2607] = 0.0;
scaleFactors[2606] = 0.0;
scaleFactors[2605] = 0.0;
scaleFactors[2604] = 0.0;
scaleFactors[2603] = 0.0;
scaleFactors[2602] = 0.0;
scaleFactors[2601] = 0.0;
scaleFactors[2600] = 0.0;
scaleFactors[2599] = 0.0;
scaleFactors[2598] = 0.0;
scaleFactors[2597] = 0.0;
scaleFactors[2596] = 0.0;
scaleFactors[2595] = 0.0;
scaleFactors[2594] = 0.0;
scaleFactors[2593] = 0.0;
scaleFactors[2592] = 0.0;
scaleFactors[2591] = 0.0;
scaleFactors[2590] = 0.0;
scaleFactors[2589] = 0.0;
scaleFactors[2588] = 0.0;
scaleFactors[2587] = 0.0;
scaleFactors[2586] = 0.0;
scaleFactors[2585] = 0.0;
scaleFactors[2584] = 0.0;
scaleFactors[2583] = 0.0;
scaleFactors[2582] = 0.0;
scaleFactors[2581] = 0.0;
scaleFactors[2580] = 0.0;
scaleFactors[2579] = 0.0;
scaleFactors[2578] = 0.0;
scaleFactors[2577] = 0.0;
scaleFactors[2576] = 0.0;
scaleFactors[2575] = 0.0;
scaleFactors[2574] = 0.0;
scaleFactors[2573] = 0.0;
scaleFactors[2572] = 0.0;
scaleFactors[2571] = 0.0;
scaleFactors[2570] = 0.0;
scaleFactors[2569] = 0.0;
scaleFactors[2568] = 0.0;
scaleFactors[2567] = 0.0;
scaleFactors[2566] = 0.0;
scaleFactors[2565] = 0.0;
scaleFactors[2564] = 0.0;
scaleFactors[2563] = 0.0;
scaleFactors[2562] = 0.0;
scaleFactors[2561] = 0.0;
scaleFactors[2560] = 0.0;
scaleFactors[2559] = 0.0;
scaleFactors[2558] = 0.0;
scaleFactors[2557] = 0.0;
scaleFactors[2556] = 0.0;
scaleFactors[2555] = 0.0;
scaleFactors[2554] = 0.0;
scaleFactors[2553] = 0.0;
scaleFactors[2552] = 0.0;
scaleFactors[2551] = 0.0;
scaleFactors[2550] = 0.0;
scaleFactors[2549] = 0.0;
scaleFactors[2548] = 0.0;
scaleFactors[2547] = 0.0;
scaleFactors[2546] = 0.0;
scaleFactors[2545] = 0.0;
scaleFactors[2544] = 0.0;
scaleFactors[2543] = 0.0;
scaleFactors[2542] = 0.0;
scaleFactors[2541] = 0.0;
scaleFactors[2540] = 0.0;
scaleFactors[2539] = 0.0;
scaleFactors[2538] = 0.0;
scaleFactors[2537] = 0.0;
scaleFactors[2536] = 0.0;
scaleFactors[2535] = 0.0;
scaleFactors[2534] = 0.0;
scaleFactors[2533] = 0.0;
scaleFactors[2532] = 0.0;
scaleFactors[2531] = 0.0;
scaleFactors[2530] = 0.0;
scaleFactors[2529] = 0.0;
scaleFactors[2528] = 0.0;
scaleFactors[2527] = 0.0;
scaleFactors[2526] = 0.0;
scaleFactors[2525] = 0.0;
scaleFactors[2524] = 0.0;
scaleFactors[2523] = 0.0;
scaleFactors[2522] = 0.0;
scaleFactors[2521] = 0.0;
scaleFactors[2520] = 0.0;
scaleFactors[2519] = 0.0;
scaleFactors[2518] = 0.0;
scaleFactors[2517] = 0.0;
scaleFactors[2516] = 0.0;
scaleFactors[2515] = 0.0;
scaleFactors[2514] = 0.0;
scaleFactors[2513] = 0.0;
scaleFactors[2512] = 0.0;
scaleFactors[2511] = 0.0;
scaleFactors[2510] = 0.0;
scaleFactors[2509] = 0.0;
scaleFactors[2508] = 0.0;
scaleFactors[2507] = 0.0;
scaleFactors[2506] = 0.0;
scaleFactors[2505] = 0.0;
scaleFactors[2504] = 0.0;
scaleFactors[2503] = 0.0;
scaleFactors[2502] = 0.0;
scaleFactors[2501] = 0.0;
scaleFactors[2500] = 0.0;
scaleFactors[2499] = 0.0;
scaleFactors[2498] = 0.0;
scaleFactors[2497] = 0.0;
scaleFactors[2496] = 0.0;
scaleFactors[2495] = 0.0;
scaleFactors[2494] = 0.0;
scaleFactors[2493] = 0.0;
scaleFactors[2492] = 0.0;
scaleFactors[2491] = 0.0;
scaleFactors[2490] = 0.0;
scaleFactors[2489] = 0.0;
scaleFactors[2488] = 0.0;
scaleFactors[2487] = 0.0;
scaleFactors[2486] = 0.0;
scaleFactors[2485] = 0.0;
scaleFactors[2484] = 0.0;
scaleFactors[2483] = 0.0;
scaleFactors[2482] = 0.0;
scaleFactors[2481] = 0.0;
scaleFactors[2480] = 0.0;
scaleFactors[2479] = 0.0;
scaleFactors[2478] = 0.0;
scaleFactors[2477] = 0.0;
scaleFactors[2476] = 0.0;
scaleFactors[2475] = 0.0;
scaleFactors[2474] = 0.0;
scaleFactors[2473] = 0.0;
scaleFactors[2472] = 0.0;
scaleFactors[2471] = 0.0;
scaleFactors[2470] = 0.0;
scaleFactors[2469] = 0.0;
scaleFactors[2468] = 0.0;
scaleFactors[2467] = 0.0;
scaleFactors[2466] = 0.0;
scaleFactors[2465] = 0.0;
scaleFactors[2464] = 0.0;
scaleFactors[2463] = 0.0;
scaleFactors[2462] = 0.0;
scaleFactors[2461] = 0.0;
scaleFactors[2460] = 0.0;
scaleFactors[2459] = 0.0;
scaleFactors[2458] = 0.0;
scaleFactors[2457] = 0.0;
scaleFactors[2456] = 0.0;
scaleFactors[2455] = 0.0;
scaleFactors[2454] = 0.0;
scaleFactors[2453] = 0.0;
scaleFactors[2452] = 0.0;
scaleFactors[2451] = 0.0;
scaleFactors[2450] = 0.0;
scaleFactors[2449] = 0.0;
scaleFactors[2448] = 0.0;
scaleFactors[2447] = 0.0;
scaleFactors[2446] = 0.0;
scaleFactors[2445] = 0.0;
scaleFactors[2444] = 0.0;
scaleFactors[2443] = 0.0;
scaleFactors[2442] = 0.0;
scaleFactors[2441] = 0.0;
scaleFactors[2440] = 0.0;
scaleFactors[2439] = 0.0;
scaleFactors[2438] = 0.0;
scaleFactors[2437] = 0.0;
scaleFactors[2436] = 0.0;
scaleFactors[2435] = 0.0;
scaleFactors[2434] = 0.0;
scaleFactors[2433] = 0.0;
scaleFactors[2432] = 0.0;
scaleFactors[2431] = 0.0;
scaleFactors[2430] = 0.0;
scaleFactors[2429] = 0.0;
scaleFactors[2428] = 0.0;
scaleFactors[2427] = 0.0;
scaleFactors[2426] = 0.0;
scaleFactors[2425] = 0.0;
scaleFactors[2424] = 0.0;
scaleFactors[2423] = 0.0;
scaleFactors[2422] = 0.0;
scaleFactors[2421] = 0.0;
scaleFactors[2420] = 0.0;
scaleFactors[2419] = 0.0;
scaleFactors[2418] = 0.0;
scaleFactors[2417] = 0.0;
scaleFactors[2416] = 0.0;
scaleFactors[2415] = 0.0;
scaleFactors[2414] = 0.0;
scaleFactors[2413] = 0.0;
scaleFactors[2412] = 0.0;
scaleFactors[2411] = 0.0;
scaleFactors[2410] = 0.0;
scaleFactors[2409] = 0.0;
scaleFactors[2408] = 0.0;
scaleFactors[2407] = 0.0;
scaleFactors[2406] = 0.0;
scaleFactors[2405] = 0.0;
scaleFactors[2404] = 0.0;
scaleFactors[2403] = 0.0;
scaleFactors[2402] = 0.0;
scaleFactors[2401] = 0.0;
scaleFactors[2400] = 0.0;
scaleFactors[2399] = 0.0;
scaleFactors[2398] = 0.0;
scaleFactors[2397] = 0.0;
scaleFactors[2396] = 0.0;
scaleFactors[2395] = 0.0;
scaleFactors[2394] = 0.0;
scaleFactors[2393] = 0.0;
scaleFactors[2392] = 0.0;
scaleFactors[2391] = 0.0;
scaleFactors[2390] = 0.0;
scaleFactors[2389] = 0.0;
scaleFactors[2388] = 0.0;
scaleFactors[2387] = 0.0;
scaleFactors[2386] = 0.0;
scaleFactors[2385] = 0.0;
scaleFactors[2384] = 0.0;
scaleFactors[2383] = 0.0;
scaleFactors[2382] = 0.0;
scaleFactors[2381] = 0.0;
scaleFactors[2380] = 0.0;
scaleFactors[2379] = 0.0;
scaleFactors[2378] = 0.0;
scaleFactors[2377] = 0.0;
scaleFactors[2376] = 0.0;
scaleFactors[2375] = 0.0;
scaleFactors[2374] = 0.0;
scaleFactors[2373] = 0.0;
scaleFactors[2372] = 0.0;
scaleFactors[2371] = 0.0;
scaleFactors[2370] = 0.0;
scaleFactors[2369] = 0.0;
scaleFactors[2368] = 0.0;
scaleFactors[2367] = 0.0;
scaleFactors[2366] = 0.0;
scaleFactors[2365] = 0.0;
scaleFactors[2364] = 0.0;
scaleFactors[2363] = 0.0;
scaleFactors[2362] = 0.0;
scaleFactors[2361] = 0.0;
scaleFactors[2360] = 0.0;
scaleFactors[2359] = 0.0;
scaleFactors[2358] = 0.0;
scaleFactors[2357] = 0.0;
scaleFactors[2356] = 0.0;
scaleFactors[2355] = 0.0;
scaleFactors[2354] = 0.0;
scaleFactors[2353] = 0.0;
scaleFactors[2352] = 0.0;
scaleFactors[2351] = 0.0;
scaleFactors[2350] = 0.0;
scaleFactors[2349] = 0.0;
scaleFactors[2348] = 0.0;
scaleFactors[2347] = 0.0;
scaleFactors[2346] = 0.0;
scaleFactors[2345] = 0.0;
scaleFactors[2344] = 0.0;
scaleFactors[2343] = 0.0;
scaleFactors[2342] = 0.0;
scaleFactors[2341] = 0.0;
scaleFactors[2340] = 0.0;
scaleFactors[2339] = 0.0;
scaleFactors[2338] = 0.0;
scaleFactors[2337] = 0.0;
scaleFactors[2336] = 0.0;
scaleFactors[2335] = 0.0;
scaleFactors[2334] = 0.0;
scaleFactors[2333] = 0.0;
scaleFactors[2332] = 0.0;
scaleFactors[2331] = 0.0;
scaleFactors[2330] = 0.0;
scaleFactors[2329] = 0.0;
scaleFactors[2328] = 0.0;
scaleFactors[2327] = 0.0;
scaleFactors[2326] = 0.0;
scaleFactors[2325] = 0.0;
scaleFactors[2324] = 0.0;
scaleFactors[2323] = 0.0;
scaleFactors[2322] = 0.0;
scaleFactors[2321] = 0.0;
scaleFactors[2320] = 0.0;
scaleFactors[2319] = 0.0;
scaleFactors[2318] = 0.0;
scaleFactors[2317] = 0.0;
scaleFactors[2316] = 0.0;
scaleFactors[2315] = 0.0;
scaleFactors[2314] = 0.0;
scaleFactors[2313] = 0.0;
scaleFactors[2312] = 0.0;
scaleFactors[2311] = 0.0;
scaleFactors[2310] = 0.0;
scaleFactors[2309] = 0.0;
scaleFactors[2308] = 0.0;
scaleFactors[2307] = 0.0;
scaleFactors[2306] = 0.0;
scaleFactors[2305] = 0.0;
scaleFactors[2304] = 0.0;
scaleFactors[2303] = 0.0;
scaleFactors[2302] = 0.0;
scaleFactors[2301] = 0.0;
scaleFactors[2300] = 0.0;
scaleFactors[2299] = 0.0;
scaleFactors[2298] = 0.0;
scaleFactors[2297] = 0.0;
scaleFactors[2296] = 0.0;
scaleFactors[2295] = 0.0;
scaleFactors[2294] = 0.0;
scaleFactors[2293] = 0.0;
scaleFactors[2292] = 0.0;
scaleFactors[2291] = 0.0;
scaleFactors[2290] = 0.0;
scaleFactors[2289] = 0.0;
scaleFactors[2288] = 0.0;
scaleFactors[2287] = 0.0;
scaleFactors[2286] = 0.0;
scaleFactors[2285] = 0.0;
scaleFactors[2284] = 0.0;
scaleFactors[2283] = 0.0;
scaleFactors[2282] = 0.0;
scaleFactors[2281] = 0.0;
scaleFactors[2280] = 0.0;
scaleFactors[2279] = 0.0;
scaleFactors[2278] = 0.0;
scaleFactors[2277] = 0.0;
scaleFactors[2276] = 0.0;
scaleFactors[2275] = 0.0;
scaleFactors[2274] = 0.0;
scaleFactors[2273] = 0.0;
scaleFactors[2272] = 0.0;
scaleFactors[2271] = 0.0;
scaleFactors[2270] = 0.0;
scaleFactors[2269] = 0.0;
scaleFactors[2268] = 0.0;
scaleFactors[2267] = 0.0;
scaleFactors[2266] = 0.0;
scaleFactors[2265] = 0.0;
scaleFactors[2264] = 0.0;
scaleFactors[2263] = 0.0;
scaleFactors[2262] = 0.0;
scaleFactors[2261] = 0.0;
scaleFactors[2260] = 0.0;
scaleFactors[2259] = 0.0;
scaleFactors[2258] = 0.0;
scaleFactors[2257] = 0.0;
scaleFactors[2256] = 0.0;
scaleFactors[2255] = 0.0;
scaleFactors[2254] = 0.0;
scaleFactors[2253] = 0.0;
scaleFactors[2252] = 0.0;
scaleFactors[2251] = 0.0;
scaleFactors[2250] = 0.0;
scaleFactors[2249] = 0.0;
scaleFactors[2248] = 0.0;
scaleFactors[2247] = 0.0;
scaleFactors[2246] = 0.0;
scaleFactors[2245] = 0.0;
scaleFactors[2244] = 0.0;
scaleFactors[2243] = 0.0;
scaleFactors[2242] = 0.0;
scaleFactors[2241] = 0.0;
scaleFactors[2240] = 0.0;
scaleFactors[2239] = 0.0;
scaleFactors[2238] = 0.0;
scaleFactors[2237] = 0.0;
scaleFactors[2236] = 0.0;
scaleFactors[2235] = 0.0;
scaleFactors[2234] = 0.0;
scaleFactors[2233] = 0.0;
scaleFactors[2232] = 0.0;
scaleFactors[2231] = 0.0;
scaleFactors[2230] = 0.0;
scaleFactors[2229] = 0.0;
scaleFactors[2228] = 0.0;
scaleFactors[2227] = 0.0;
scaleFactors[2226] = 0.0;
scaleFactors[2225] = 0.0;
scaleFactors[2224] = 0.0;
scaleFactors[2223] = 0.0;
scaleFactors[2222] = 0.0;
scaleFactors[2221] = 0.0;
scaleFactors[2220] = 0.0;
scaleFactors[2219] = 0.0;
scaleFactors[2218] = 0.0;
scaleFactors[2217] = 0.0;
scaleFactors[2216] = 0.0;
scaleFactors[2215] = 0.0;
scaleFactors[2214] = 0.0;
scaleFactors[2213] = 0.0;
scaleFactors[2212] = 0.0;
scaleFactors[2211] = 0.0;
scaleFactors[2210] = 0.0;
scaleFactors[2209] = 0.0;
scaleFactors[2208] = 0.0;
scaleFactors[2207] = 0.0;
scaleFactors[2206] = 0.0;
scaleFactors[2205] = 0.0;
scaleFactors[2204] = 0.0;
scaleFactors[2203] = 0.0;
scaleFactors[2202] = 0.0;
scaleFactors[2201] = 0.0;
scaleFactors[2200] = 0.0;
scaleFactors[2199] = 0.0;
scaleFactors[2198] = 0.0;
scaleFactors[2197] = 0.0;
scaleFactors[2196] = 0.0;
scaleFactors[2195] = 0.0;
scaleFactors[2194] = 0.0;
scaleFactors[2193] = 0.0;
scaleFactors[2192] = 0.0;
scaleFactors[2191] = 0.0;
scaleFactors[2190] = 0.0;
scaleFactors[2189] = 0.0;
scaleFactors[2188] = 0.0;
scaleFactors[2187] = 0.0;
scaleFactors[2186] = 0.0;
scaleFactors[2185] = 0.0;
scaleFactors[2184] = 0.0;
scaleFactors[2183] = 0.0;
scaleFactors[2182] = 0.0;
scaleFactors[2181] = 0.0;
scaleFactors[2180] = 0.0;
scaleFactors[2179] = 0.0;
scaleFactors[2178] = 0.0;
scaleFactors[2177] = 0.0;
scaleFactors[2176] = 0.0;
scaleFactors[2175] = 0.0;
scaleFactors[2174] = 0.0;
scaleFactors[2173] = 0.0;
scaleFactors[2172] = 0.0;
scaleFactors[2171] = 0.0;
scaleFactors[2170] = 0.0;
scaleFactors[2169] = 0.0;
scaleFactors[2168] = 0.0;
scaleFactors[2167] = 0.0;
scaleFactors[2166] = 0.0;
scaleFactors[2165] = 0.0;
scaleFactors[2164] = 0.0;
scaleFactors[2163] = 0.0;
scaleFactors[2162] = 0.0;
scaleFactors[2161] = 0.0;
scaleFactors[2160] = 0.0;
scaleFactors[2159] = 0.0;
scaleFactors[2158] = 0.0;
scaleFactors[2157] = 0.0;
scaleFactors[2156] = 0.0;
scaleFactors[2155] = 0.0;
scaleFactors[2154] = 0.0;
scaleFactors[2153] = 0.0;
scaleFactors[2152] = 0.0;
scaleFactors[2151] = 0.0;
scaleFactors[2150] = 0.0;
scaleFactors[2149] = 0.0;
scaleFactors[2148] = 0.0;
scaleFactors[2147] = 0.0;
scaleFactors[2146] = 0.0;
scaleFactors[2145] = 0.0;
scaleFactors[2144] = 0.0;
scaleFactors[2143] = 0.0;
scaleFactors[2142] = 0.0;
scaleFactors[2141] = 0.0;
scaleFactors[2140] = 0.0;
scaleFactors[2139] = 0.0;
scaleFactors[2138] = 0.0;
scaleFactors[2137] = 0.0;
scaleFactors[2136] = 0.0;
scaleFactors[2135] = 0.0;
scaleFactors[2134] = 0.0;
scaleFactors[2133] = 0.0;
scaleFactors[2132] = 0.0;
scaleFactors[2131] = 0.0;
scaleFactors[2130] = 0.0;
scaleFactors[2129] = 0.0;
scaleFactors[2128] = 0.0;
scaleFactors[2127] = 0.0;
scaleFactors[2126] = 0.0;
scaleFactors[2125] = 0.0;
scaleFactors[2124] = 0.0;
scaleFactors[2123] = 0.0;
scaleFactors[2122] = 0.0;
scaleFactors[2121] = 0.0;
scaleFactors[2120] = 0.0;
scaleFactors[2119] = 0.0;
scaleFactors[2118] = 0.0;
scaleFactors[2117] = 0.0;
scaleFactors[2116] = 0.0;
scaleFactors[2115] = 0.0;
scaleFactors[2114] = 0.0;
scaleFactors[2113] = 0.0;
scaleFactors[2112] = 0.0;
scaleFactors[2111] = 0.0;
scaleFactors[2110] = 0.0;
scaleFactors[2109] = 0.0;
scaleFactors[2108] = 0.0;
scaleFactors[2107] = 0.0;
scaleFactors[2106] = 0.0;
scaleFactors[2105] = 0.0;
scaleFactors[2104] = 0.0;
scaleFactors[2103] = 0.0;
scaleFactors[2102] = 0.0;
scaleFactors[2101] = 0.0;
scaleFactors[2100] = 0.0;
scaleFactors[2099] = 0.0;
scaleFactors[2098] = 0.0;
scaleFactors[2097] = 0.0;
scaleFactors[2096] = 0.0;
scaleFactors[2095] = 0.0;
scaleFactors[2094] = 0.0;
scaleFactors[2093] = 0.0;
scaleFactors[2092] = 0.0;
scaleFactors[2091] = 0.0;
scaleFactors[2090] = 0.0;
scaleFactors[2089] = 0.0;
scaleFactors[2088] = 0.0;
scaleFactors[2087] = 0.0;
scaleFactors[2086] = 0.0;
scaleFactors[2085] = 0.0;
scaleFactors[2084] = 0.0;
scaleFactors[2083] = 0.0;
scaleFactors[2082] = 0.0;
scaleFactors[2081] = 0.0;
scaleFactors[2080] = 0.0;
scaleFactors[2079] = 0.0;
scaleFactors[2078] = 0.0;
scaleFactors[2077] = 0.0;
scaleFactors[2076] = 0.0;
scaleFactors[2075] = 0.0;
scaleFactors[2074] = 0.0;
scaleFactors[2073] = 0.0;
scaleFactors[2072] = 0.0;
scaleFactors[2071] = 0.0;
scaleFactors[2070] = 0.0;
scaleFactors[2069] = 0.0;
scaleFactors[2068] = 0.0;
scaleFactors[2067] = 0.0;
scaleFactors[2066] = 0.0;
scaleFactors[2065] = 0.0;
scaleFactors[2064] = 0.0;
scaleFactors[2063] = 0.0;
scaleFactors[2062] = 0.0;
scaleFactors[2061] = 0.0;
scaleFactors[2060] = 0.0;
scaleFactors[2059] = 0.0;
scaleFactors[2058] = 0.0;
scaleFactors[2057] = 0.0;
scaleFactors[2056] = 0.0;
scaleFactors[2055] = 0.0;
scaleFactors[2054] = 0.0;
scaleFactors[2053] = 0.0;
scaleFactors[2052] = 0.0;
scaleFactors[2051] = 0.0;
scaleFactors[2050] = 0.0;
scaleFactors[2049] = 0.0;
scaleFactors[2048] = 0.0;
scaleFactors[2047] = 0.0;
scaleFactors[2046] = 0.0;
scaleFactors[2045] = 0.0;
scaleFactors[2044] = 0.0;
scaleFactors[2043] = 0.0;
scaleFactors[2042] = 0.0;
scaleFactors[2041] = 0.0;
scaleFactors[2040] = 0.0;
scaleFactors[2039] = 0.0;
scaleFactors[2038] = 0.0;
scaleFactors[2037] = 0.0;
scaleFactors[2036] = 0.0;
scaleFactors[2035] = 0.0;
scaleFactors[2034] = 0.0;
scaleFactors[2033] = 0.0;
scaleFactors[2032] = 0.0;
scaleFactors[2031] = 0.0;
scaleFactors[2030] = 0.0;
scaleFactors[2029] = 0.0;
scaleFactors[2028] = 0.0;
scaleFactors[2027] = 0.0;
scaleFactors[2026] = 0.0;
scaleFactors[2025] = 0.0;
scaleFactors[2024] = 0.0;
scaleFactors[2023] = 0.0;
scaleFactors[2022] = 0.0;
scaleFactors[2021] = 0.0;
scaleFactors[2020] = 0.0;
scaleFactors[2019] = 0.0;
scaleFactors[2018] = 0.0;
scaleFactors[2017] = 0.0;
scaleFactors[2016] = 0.0;
scaleFactors[2015] = 0.0;
scaleFactors[2014] = 0.0;
scaleFactors[2013] = 0.0;
scaleFactors[2012] = 0.0;
scaleFactors[2011] = 0.0;
scaleFactors[2010] = 0.0;
scaleFactors[2009] = 0.0;
scaleFactors[2008] = 0.0;
scaleFactors[2007] = 0.0;
scaleFactors[2006] = 0.0;
scaleFactors[2005] = 0.0;
scaleFactors[2004] = 0.0;
scaleFactors[2003] = 0.0;
scaleFactors[2002] = 0.0;
scaleFactors[2001] = 0.0;
scaleFactors[2000] = 0.0;
scaleFactors[1999] = 0.0;
scaleFactors[1998] = 0.0;
scaleFactors[1997] = 0.0;
scaleFactors[1996] = 0.0;
scaleFactors[1995] = 0.0;
scaleFactors[1994] = 0.0;
scaleFactors[1993] = 0.0;
scaleFactors[1992] = 0.0;
scaleFactors[1991] = 0.0;
scaleFactors[1990] = 0.0;
scaleFactors[1989] = 0.0;
scaleFactors[1988] = 0.0;
scaleFactors[1987] = 0.0;
scaleFactors[1986] = 0.0;
scaleFactors[1985] = 0.0;
scaleFactors[1984] = 0.0;
scaleFactors[1983] = 0.0;
scaleFactors[1982] = 0.0;
scaleFactors[1981] = 0.0;
scaleFactors[1980] = 0.0;
scaleFactors[1979] = 0.0;
scaleFactors[1978] = 0.0;
scaleFactors[1977] = 0.0;
scaleFactors[1976] = 0.0;
scaleFactors[1975] = 0.0;
scaleFactors[1974] = 0.0;
scaleFactors[1973] = 0.0;
scaleFactors[1972] = 0.0;
scaleFactors[1971] = 0.0;
scaleFactors[1970] = 0.0;
scaleFactors[1969] = 0.0;
scaleFactors[1968] = 0.0;
scaleFactors[1967] = 0.0;
scaleFactors[1966] = 0.0;
scaleFactors[1965] = 0.0;
scaleFactors[1964] = 0.0;
scaleFactors[1963] = 0.0;
scaleFactors[1962] = 0.0;
scaleFactors[1961] = 0.0;
scaleFactors[1960] = 0.0;
scaleFactors[1959] = 0.0;
scaleFactors[1958] = 0.0;
scaleFactors[1957] = 0.0;
scaleFactors[1956] = 0.0;
scaleFactors[1955] = 0.0;
scaleFactors[1954] = 0.0;
scaleFactors[1953] = 0.0;
scaleFactors[1952] = 0.0;
scaleFactors[1951] = 0.0;
scaleFactors[1950] = 0.0;
scaleFactors[1949] = 0.0;
scaleFactors[1948] = 0.0;
scaleFactors[1947] = 0.0;
scaleFactors[1946] = 0.0;
scaleFactors[1945] = 0.0;
scaleFactors[1944] = 0.0;
scaleFactors[1943] = 0.0;
scaleFactors[1942] = 0.0;
scaleFactors[1941] = 0.0;
scaleFactors[1940] = 0.0;
scaleFactors[1939] = 0.0;
scaleFactors[1938] = 0.0;
scaleFactors[1937] = 0.0;
scaleFactors[1936] = 0.0;
scaleFactors[1935] = 0.0;
scaleFactors[1934] = 0.0;
scaleFactors[1933] = 0.0;
scaleFactors[1932] = 0.0;
scaleFactors[1931] = 0.0;
scaleFactors[1930] = 0.0;
scaleFactors[1929] = 0.0;
scaleFactors[1928] = 0.0;
scaleFactors[1927] = 0.0;
scaleFactors[1926] = 0.0;
scaleFactors[1925] = 0.0;
scaleFactors[1924] = 0.0;
scaleFactors[1923] = 0.0;
scaleFactors[1922] = 0.0;
scaleFactors[1921] = 0.0;
scaleFactors[1920] = 0.0;
scaleFactors[1919] = 0.0;
scaleFactors[1918] = 0.0;
scaleFactors[1917] = 0.0;
scaleFactors[1916] = 0.0;
scaleFactors[1915] = 0.0;
scaleFactors[1914] = 0.0;
scaleFactors[1913] = 0.0;
scaleFactors[1912] = 0.0;
scaleFactors[1911] = 0.0;
scaleFactors[1910] = 0.0;
scaleFactors[1909] = 0.0;
scaleFactors[1908] = 0.0;
scaleFactors[1907] = 0.0;
scaleFactors[1906] = 0.0;
scaleFactors[1905] = 0.0;
scaleFactors[1904] = 0.0;
scaleFactors[1903] = 0.0;
scaleFactors[1902] = 0.0;
scaleFactors[1901] = 0.0;
scaleFactors[1900] = 0.0;
scaleFactors[1899] = 0.0;
scaleFactors[1898] = 0.0;
scaleFactors[1897] = 0.0;
scaleFactors[1896] = 0.0;
scaleFactors[1895] = 0.0;
scaleFactors[1894] = 0.0;
scaleFactors[1893] = 0.0;
scaleFactors[1892] = 0.0;
scaleFactors[1891] = 0.0;
scaleFactors[1890] = 0.0;
scaleFactors[1889] = 0.0;
scaleFactors[1888] = 0.0;
scaleFactors[1887] = 0.0;
scaleFactors[1886] = 0.0;
scaleFactors[1885] = 0.0;
scaleFactors[1884] = 0.0;
scaleFactors[1883] = 0.0;
scaleFactors[1882] = 0.0;
scaleFactors[1881] = 0.0;
scaleFactors[1880] = 0.0;
scaleFactors[1879] = 0.0;
scaleFactors[1878] = 0.0;
scaleFactors[1877] = 0.0;
scaleFactors[1876] = 0.0;
scaleFactors[1875] = 0.0;
scaleFactors[1874] = 0.0;
scaleFactors[1873] = 0.0;
scaleFactors[1872] = 0.0;
scaleFactors[1871] = 0.0;
scaleFactors[1870] = 0.0;
scaleFactors[1869] = 0.0;
scaleFactors[1868] = 0.0;
scaleFactors[1867] = 0.0;
scaleFactors[1866] = 0.0;
scaleFactors[1865] = 0.0;
scaleFactors[1864] = 0.0;
scaleFactors[1863] = 0.0;
scaleFactors[1862] = 0.0;
scaleFactors[1861] = 0.0;
scaleFactors[1860] = 0.0;
scaleFactors[1859] = 0.0;
scaleFactors[1858] = 0.0;
scaleFactors[1857] = 0.0;
scaleFactors[1856] = 0.0;
scaleFactors[1855] = 0.0;
scaleFactors[1854] = 0.0;
scaleFactors[1853] = 0.0;
scaleFactors[1852] = 0.0;
scaleFactors[1851] = 0.0;
scaleFactors[1850] = 0.0;
scaleFactors[1849] = 0.0;
scaleFactors[1848] = 0.0;
scaleFactors[1847] = 0.0;
scaleFactors[1846] = 0.0;
scaleFactors[1845] = 0.0;
scaleFactors[1844] = 0.0;
scaleFactors[1843] = 0.0;
scaleFactors[1842] = 0.0;
scaleFactors[1841] = 0.0;
scaleFactors[1840] = 0.0;
scaleFactors[1839] = 0.0;
scaleFactors[1838] = 0.0;
scaleFactors[1837] = 0.0;
scaleFactors[1836] = 0.0;
scaleFactors[1835] = 0.0;
scaleFactors[1834] = 0.0;
scaleFactors[1833] = 0.0;
scaleFactors[1832] = 0.0;
scaleFactors[1831] = 0.0;
scaleFactors[1830] = 0.0;
scaleFactors[1829] = 0.0;
scaleFactors[1828] = 0.0;
scaleFactors[1827] = 0.0;
scaleFactors[1826] = 0.0;
scaleFactors[1825] = 0.0;
scaleFactors[1824] = 0.0;
scaleFactors[1823] = 0.0;
scaleFactors[1822] = 0.0;
scaleFactors[1821] = 0.0;
scaleFactors[1820] = 0.0;
scaleFactors[1819] = 0.0;
scaleFactors[1818] = 0.0;
scaleFactors[1817] = 0.0;
scaleFactors[1816] = 0.0;
scaleFactors[1815] = 0.0;
scaleFactors[1814] = 0.0;
scaleFactors[1813] = 0.0;
scaleFactors[1812] = 0.0;
scaleFactors[1811] = 0.0;
scaleFactors[1810] = 0.0;
scaleFactors[1809] = 0.0;
scaleFactors[1808] = 0.0;
scaleFactors[1807] = 0.0;
scaleFactors[1806] = 0.0;
scaleFactors[1805] = 0.0;
scaleFactors[1804] = 0.0;
scaleFactors[1803] = 0.0;
scaleFactors[1802] = 0.0;
scaleFactors[1801] = 0.0;
scaleFactors[1800] = 0.0;
scaleFactors[1799] = 0.0;
scaleFactors[1798] = 0.0;
scaleFactors[1797] = 0.0;
scaleFactors[1796] = 0.0;
scaleFactors[1795] = 0.0;
scaleFactors[1794] = 0.0;
scaleFactors[1793] = 0.0;
scaleFactors[1792] = 0.0;
scaleFactors[1791] = 0.0;
scaleFactors[1790] = 0.0;
scaleFactors[1789] = 0.0;
scaleFactors[1788] = 0.0;
scaleFactors[1787] = 0.0;
scaleFactors[1786] = 0.0;
scaleFactors[1785] = 0.0;
scaleFactors[1784] = 0.0;
scaleFactors[1783] = 0.0;
scaleFactors[1782] = 0.0;
scaleFactors[1781] = 0.0;
scaleFactors[1780] = 0.0;
scaleFactors[1779] = 0.0;
scaleFactors[1778] = 0.0;
scaleFactors[1777] = 0.0;
scaleFactors[1776] = 0.0;
scaleFactors[1775] = 0.0;
scaleFactors[1774] = 0.0;
scaleFactors[1773] = 0.0;
scaleFactors[1772] = 0.0;
scaleFactors[1771] = 0.0;
scaleFactors[1770] = 0.0;
scaleFactors[1769] = 0.0;
scaleFactors[1768] = 0.0;
scaleFactors[1767] = 0.0;
scaleFactors[1766] = 0.0;
scaleFactors[1765] = 0.0;
scaleFactors[1764] = 0.0;
scaleFactors[1763] = 0.0;
scaleFactors[1762] = 0.0;
scaleFactors[1761] = 0.0;
scaleFactors[1760] = 0.0;
scaleFactors[1759] = 0.0;
scaleFactors[1758] = 0.0;
scaleFactors[1757] = 0.0;
scaleFactors[1756] = 0.0;
scaleFactors[1755] = 0.0;
scaleFactors[1754] = 0.0;
scaleFactors[1753] = 0.0;
scaleFactors[1752] = 0.0;
scaleFactors[1751] = 0.0;
scaleFactors[1750] = 0.0;
scaleFactors[1749] = 0.0;
scaleFactors[1748] = 0.0;
scaleFactors[1747] = 0.0;
scaleFactors[1746] = 0.0;
scaleFactors[1745] = 0.0;
scaleFactors[1744] = 0.0;
scaleFactors[1743] = 0.0;
scaleFactors[1742] = 0.0;
scaleFactors[1741] = 0.0;
scaleFactors[1740] = 0.0;
scaleFactors[1739] = 0.0;
scaleFactors[1738] = 0.0;
scaleFactors[1737] = 0.0;
scaleFactors[1736] = 0.0;
scaleFactors[1735] = 0.0;
scaleFactors[1734] = 0.0;
scaleFactors[1733] = 0.0;
scaleFactors[1732] = 0.0;
scaleFactors[1731] = 0.0;
scaleFactors[1730] = 0.0;
scaleFactors[1729] = 0.0;
scaleFactors[1728] = 0.0;
scaleFactors[1727] = 0.0;
scaleFactors[1726] = 0.0;
scaleFactors[1725] = 0.0;
scaleFactors[1724] = 0.0;
scaleFactors[1723] = 0.0;
scaleFactors[1722] = 0.0;
scaleFactors[1721] = 0.0;
scaleFactors[1720] = 0.0;
scaleFactors[1719] = 0.0;
scaleFactors[1718] = 0.0;
scaleFactors[1717] = 0.0;
scaleFactors[1716] = 0.0;
scaleFactors[1715] = 0.0;
scaleFactors[1714] = 0.0;
scaleFactors[1713] = 0.0;
scaleFactors[1712] = 0.0;
scaleFactors[1711] = 0.0;
scaleFactors[1710] = 0.0;
scaleFactors[1709] = 0.0;
scaleFactors[1708] = 0.0;
scaleFactors[1707] = 0.0;
scaleFactors[1706] = 0.0;
scaleFactors[1705] = 0.0;
scaleFactors[1704] = 0.0;
scaleFactors[1703] = 0.0;
scaleFactors[1702] = 0.0;
scaleFactors[1701] = 0.0;
scaleFactors[1700] = 0.0;
scaleFactors[1699] = 0.0;
scaleFactors[1698] = 0.0;
scaleFactors[1697] = 0.0;
scaleFactors[1696] = 0.0;
scaleFactors[1695] = 0.0;
scaleFactors[1694] = 0.0;
scaleFactors[1693] = 0.0;
scaleFactors[1692] = 0.0;
scaleFactors[1691] = 0.0;
scaleFactors[1690] = 0.0;
scaleFactors[1689] = 0.0;
scaleFactors[1688] = 0.0;
scaleFactors[1687] = 0.0;
scaleFactors[1686] = 0.0;
scaleFactors[1685] = 0.0;
scaleFactors[1684] = 0.0;
scaleFactors[1683] = 0.0;
scaleFactors[1682] = 0.0;
scaleFactors[1681] = 0.0;
scaleFactors[1680] = 0.0;
scaleFactors[1679] = 0.0;
scaleFactors[1678] = 0.0;
scaleFactors[1677] = 0.0;
scaleFactors[1676] = 0.0;
scaleFactors[1675] = 0.0;
scaleFactors[1674] = 0.0;
scaleFactors[1673] = 0.0;
scaleFactors[1672] = 0.0;
scaleFactors[1671] = 0.0;
scaleFactors[1670] = 0.0;
scaleFactors[1669] = 0.0;
scaleFactors[1668] = 0.0;
scaleFactors[1667] = 0.0;
scaleFactors[1666] = 0.0;
scaleFactors[1665] = 0.0;
scaleFactors[1664] = 0.0;
scaleFactors[1663] = 0.0;
scaleFactors[1662] = 0.0;
scaleFactors[1661] = 0.0;
scaleFactors[1660] = 0.0;
scaleFactors[1659] = 0.0;
scaleFactors[1658] = 0.0;
scaleFactors[1657] = 0.0;
scaleFactors[1656] = 0.0;
scaleFactors[1655] = 0.0;
scaleFactors[1654] = 0.0;
scaleFactors[1653] = 0.0;
scaleFactors[1652] = 0.0;
scaleFactors[1651] = 0.0;
scaleFactors[1650] = 0.0;
scaleFactors[1649] = 0.0;
scaleFactors[1648] = 0.0;
scaleFactors[1647] = 0.0;
scaleFactors[1646] = 0.0;
scaleFactors[1645] = 0.0;
scaleFactors[1644] = 0.0;
scaleFactors[1643] = 0.0;
scaleFactors[1642] = 0.0;
scaleFactors[1641] = 0.0;
scaleFactors[1640] = 0.0;
scaleFactors[1639] = 0.0;
scaleFactors[1638] = 0.0;
scaleFactors[1637] = 0.0;
scaleFactors[1636] = 0.0;
scaleFactors[1635] = 0.0;
scaleFactors[1634] = 0.0;
scaleFactors[1633] = 0.0;
scaleFactors[1632] = 0.0;
scaleFactors[1631] = 0.0;
scaleFactors[1630] = 0.0;
scaleFactors[1629] = 0.0;
scaleFactors[1628] = 0.0;
scaleFactors[1627] = 0.0;
scaleFactors[1626] = 0.0;
scaleFactors[1625] = 0.0;
scaleFactors[1624] = 0.0;
scaleFactors[1623] = 0.0;
scaleFactors[1622] = 0.0;
scaleFactors[1621] = 0.0;
scaleFactors[1620] = 0.0;
scaleFactors[1619] = 0.0;
scaleFactors[1618] = 0.0;
scaleFactors[1617] = 0.0;
scaleFactors[1616] = 0.0;
scaleFactors[1615] = 0.0;
scaleFactors[1614] = 0.0;
scaleFactors[1613] = 0.0;
scaleFactors[1612] = 0.0;
scaleFactors[1611] = 0.0;
scaleFactors[1610] = 0.0;
scaleFactors[1609] = 0.0;
scaleFactors[1608] = 0.0;
scaleFactors[1607] = 0.0;
scaleFactors[1606] = 0.0;
scaleFactors[1605] = 0.0;
scaleFactors[1604] = 0.0;
scaleFactors[1603] = 0.0;
scaleFactors[1602] = 0.0;
scaleFactors[1601] = 0.0;
scaleFactors[1600] = 0.0;
scaleFactors[1599] = 0.0;
scaleFactors[1598] = 0.0;
scaleFactors[1597] = 0.0;
scaleFactors[1596] = 0.0;
scaleFactors[1595] = 0.0;
scaleFactors[1594] = 0.0;
scaleFactors[1593] = 0.0;
scaleFactors[1592] = 0.0;
scaleFactors[1591] = 0.0;
scaleFactors[1590] = 0.0;
scaleFactors[1589] = 0.0;
scaleFactors[1588] = 0.0;
scaleFactors[1587] = 0.0;
scaleFactors[1586] = 0.0;
scaleFactors[1585] = 0.0;
scaleFactors[1584] = 0.0;
scaleFactors[1583] = 0.0;
scaleFactors[1582] = 0.0;
scaleFactors[1581] = 0.0;
scaleFactors[1580] = 0.0;
scaleFactors[1579] = 0.0;
scaleFactors[1578] = 0.0;
scaleFactors[1577] = 0.0;
scaleFactors[1576] = 0.0;
scaleFactors[1575] = 0.0;
scaleFactors[1574] = 0.0;
scaleFactors[1573] = 0.0;
scaleFactors[1572] = 0.0;
scaleFactors[1571] = 0.0;
scaleFactors[1570] = 0.0;
scaleFactors[1569] = 0.0;
scaleFactors[1568] = 0.0;
scaleFactors[1567] = 0.0;
scaleFactors[1566] = 0.0;
scaleFactors[1565] = 0.0;
scaleFactors[1564] = 0.0;
scaleFactors[1563] = 0.0;
scaleFactors[1562] = 0.0;
scaleFactors[1561] = 0.0;
scaleFactors[1560] = 0.0;
scaleFactors[1559] = 0.0;
scaleFactors[1558] = 0.0;
scaleFactors[1557] = 0.0;
scaleFactors[1556] = 0.0;
scaleFactors[1555] = 0.0;
scaleFactors[1554] = 0.0;
scaleFactors[1553] = 0.0;
scaleFactors[1552] = 0.0;
scaleFactors[1551] = 0.0;
scaleFactors[1550] = 0.0;
scaleFactors[1549] = 0.0;
scaleFactors[1548] = 0.0;
scaleFactors[1547] = 0.0;
scaleFactors[1546] = 0.0;
scaleFactors[1545] = 0.0;
scaleFactors[1544] = 0.0;
scaleFactors[1543] = 0.0;
scaleFactors[1542] = 0.0;
scaleFactors[1541] = 0.0;
scaleFactors[1540] = 0.0;
scaleFactors[1539] = 0.0;
scaleFactors[1538] = 0.0;
scaleFactors[1537] = 0.0;
scaleFactors[1536] = 0.0;
scaleFactors[1535] = 0.0;
scaleFactors[1534] = 0.0;
scaleFactors[1533] = 0.0;
scaleFactors[1532] = 0.0;
scaleFactors[1531] = 0.0;
scaleFactors[1530] = 0.0;
scaleFactors[1529] = 0.0;
scaleFactors[1528] = 0.0;
scaleFactors[1527] = 0.0;
scaleFactors[1526] = 0.0;
scaleFactors[1525] = 0.0;
scaleFactors[1524] = 0.0;
scaleFactors[1523] = 0.0;
scaleFactors[1522] = 0.0;
scaleFactors[1521] = 0.0;
scaleFactors[1520] = 0.0;
scaleFactors[1519] = 0.0;
scaleFactors[1518] = 0.0;
scaleFactors[1517] = 0.0;
scaleFactors[1516] = 0.0;
scaleFactors[1515] = 0.0;
scaleFactors[1514] = 0.0;
scaleFactors[1513] = 0.0;
scaleFactors[1512] = 0.0;
scaleFactors[1511] = 0.0;
scaleFactors[1510] = 0.0;
scaleFactors[1509] = 0.0;
scaleFactors[1508] = 0.0;
scaleFactors[1507] = 0.0;
scaleFactors[1506] = 0.0;
scaleFactors[1505] = 0.0;
scaleFactors[1504] = 0.0;
scaleFactors[1503] = 0.0;
scaleFactors[1502] = 0.0;
scaleFactors[1501] = 0.0;
scaleFactors[1500] = 0.0;
scaleFactors[1499] = 0.0;
scaleFactors[1498] = 0.0;
scaleFactors[1497] = 0.0;
scaleFactors[1496] = 0.0;
scaleFactors[1495] = 0.0;
scaleFactors[1494] = 0.0;
scaleFactors[1493] = 0.0;
scaleFactors[1492] = 0.0;
scaleFactors[1491] = 0.0;
scaleFactors[1490] = 0.0;
scaleFactors[1489] = 00.000100;
scaleFactors[1488] = 00.000101;
scaleFactors[1487] = 00.000103;
scaleFactors[1486] = 00.000104;
scaleFactors[1485] = 00.000105;
scaleFactors[1484] = 00.000107;
scaleFactors[1483] = 00.000108;
scaleFactors[1482] = 00.000110;
scaleFactors[1481] = 00.000111;
scaleFactors[1480] = 00.000112;
scaleFactors[1479] = 00.000114;
scaleFactors[1478] = 00.000115;
scaleFactors[1477] = 00.000117;
scaleFactors[1476] = 00.000118;
scaleFactors[1475] = 00.000120;
scaleFactors[1474] = 00.000122;
scaleFactors[1473] = 00.000123;
scaleFactors[1472] = 00.000125;
scaleFactors[1471] = 00.000126;
scaleFactors[1470] = 00.000128;
scaleFactors[1469] = 00.000130;
scaleFactors[1468] = 00.000131;
scaleFactors[1467] = 00.000133;
scaleFactors[1466] = 00.000135;
scaleFactors[1465] = 00.000137;
scaleFactors[1464] = 00.000138;
scaleFactors[1463] = 00.000140;
scaleFactors[1462] = 00.000142;
scaleFactors[1461] = 00.000144;
scaleFactors[1460] = 00.000146;
scaleFactors[1459] = 00.000148;
scaleFactors[1458] = 00.000150;
scaleFactors[1457] = 00.000152;
scaleFactors[1456] = 00.000154;
scaleFactors[1455] = 00.000156;
scaleFactors[1454] = 00.000158;
scaleFactors[1453] = 00.000160;
scaleFactors[1452] = 00.000162;
scaleFactors[1451] = 00.000164;
scaleFactors[1450] = 00.000166;
scaleFactors[1449] = 00.000168;
scaleFactors[1448] = 00.000171;
scaleFactors[1447] = 00.000173;
scaleFactors[1446] = 00.000175;
scaleFactors[1445] = 00.000177;
scaleFactors[1444] = 00.000180;
scaleFactors[1443] = 00.000182;
scaleFactors[1442] = 00.000184;
scaleFactors[1441] = 00.000187;
scaleFactors[1440] = 00.000189;
scaleFactors[1439] = 00.000192;
scaleFactors[1438] = 00.000194;
scaleFactors[1437] = 00.000197;
scaleFactors[1436] = 00.000199;
scaleFactors[1435] = 00.000202;
scaleFactors[1434] = 00.000205;
scaleFactors[1433] = 00.000207;
scaleFactors[1432] = 00.000210;
scaleFactors[1431] = 00.000213;
scaleFactors[1430] = 00.000216;
scaleFactors[1429] = 00.000218;
scaleFactors[1428] = 00.000221;
scaleFactors[1427] = 00.000224;
scaleFactors[1426] = 00.000227;
scaleFactors[1425] = 00.000230;
scaleFactors[1424] = 00.000233;
scaleFactors[1423] = 00.000236;
scaleFactors[1422] = 00.000239;
scaleFactors[1421] = 00.000242;
scaleFactors[1420] = 00.000245;
scaleFactors[1419] = 00.000249;
scaleFactors[1418] = 00.000252;
scaleFactors[1417] = 00.000255;
scaleFactors[1416] = 00.000259;
scaleFactors[1415] = 00.000262;
scaleFactors[1414] = 00.000265;
scaleFactors[1413] = 00.000269;
scaleFactors[1412] = 00.000272;
scaleFactors[1411] = 00.000276;
scaleFactors[1410] = 00.000280;
scaleFactors[1409] = 00.000283;
scaleFactors[1408] = 00.000287;
scaleFactors[1407] = 00.000291;
scaleFactors[1406] = 00.000295;
scaleFactors[1405] = 00.000298;
scaleFactors[1404] = 00.000302;
scaleFactors[1403] = 00.000306;
scaleFactors[1402] = 00.000310;
scaleFactors[1401] = 00.000314;
scaleFactors[1400] = 00.000318;
scaleFactors[1399] = 00.000323;
scaleFactors[1398] = 00.000327;
scaleFactors[1397] = 00.000331;
scaleFactors[1396] = 00.000335;
scaleFactors[1395] = 00.000340;
scaleFactors[1394] = 00.000344;
scaleFactors[1393] = 00.000349;
scaleFactors[1392] = 00.000353;
scaleFactors[1391] = 00.000358;
scaleFactors[1390] = 00.000363;
scaleFactors[1389] = 00.000367;
scaleFactors[1388] = 00.000372;
scaleFactors[1387] = 00.000377;
scaleFactors[1386] = 00.000382;
scaleFactors[1385] = 00.000387;
scaleFactors[1384] = 00.000392;
scaleFactors[1383] = 00.000397;
scaleFactors[1382] = 00.000403;
scaleFactors[1381] = 00.000408;
scaleFactors[1380] = 00.000413;
scaleFactors[1379] = 00.000419;
scaleFactors[1378] = 00.000424;
scaleFactors[1377] = 00.000430;
scaleFactors[1376] = 00.000435;
scaleFactors[1375] = 00.000441;
scaleFactors[1374] = 00.000447;
scaleFactors[1373] = 00.000453;
scaleFactors[1372] = 00.000458;
scaleFactors[1371] = 00.000464;
scaleFactors[1370] = 00.000471;
scaleFactors[1369] = 00.000477;
scaleFactors[1368] = 00.000483;
scaleFactors[1367] = 00.000489;
scaleFactors[1366] = 00.000496;
scaleFactors[1365] = 00.000502;
scaleFactors[1364] = 00.000509;
scaleFactors[1363] = 00.000515;
scaleFactors[1362] = 00.000522;
scaleFactors[1361] = 00.000529;
scaleFactors[1360] = 00.000536;
scaleFactors[1359] = 00.000543;
scaleFactors[1358] = 00.000550;
scaleFactors[1357] = 00.000557;
scaleFactors[1356] = 00.000565;
scaleFactors[1355] = 00.000572;
scaleFactors[1354] = 00.000580;
scaleFactors[1353] = 00.000587;
scaleFactors[1352] = 00.000595;
scaleFactors[1351] = 00.000603;
scaleFactors[1350] = 00.000610;
scaleFactors[1349] = 00.000618;
scaleFactors[1348] = 00.000627;
scaleFactors[1347] = 00.000635;
scaleFactors[1346] = 00.000643;
scaleFactors[1345] = 00.000652;
scaleFactors[1344] = 00.000660;
scaleFactors[1343] = 00.000669;
scaleFactors[1342] = 00.000677;
scaleFactors[1341] = 00.000686;
scaleFactors[1340] = 00.000695;
scaleFactors[1339] = 00.000704;
scaleFactors[1338] = 00.000714;
scaleFactors[1337] = 00.000723;
scaleFactors[1336] = 00.000732;
scaleFactors[1335] = 00.000742;
scaleFactors[1334] = 00.000752;
scaleFactors[1333] = 00.000762;
scaleFactors[1332] = 00.000772;
scaleFactors[1331] = 00.000782;
scaleFactors[1330] = 00.000792;
scaleFactors[1329] = 00.000802;
scaleFactors[1328] = 00.000813;
scaleFactors[1327] = 00.000824;
scaleFactors[1326] = 00.000834;
scaleFactors[1325] = 00.000845;
scaleFactors[1324] = 00.000856;
scaleFactors[1323] = 00.000868;
scaleFactors[1322] = 00.000879;
scaleFactors[1321] = 00.000890;
scaleFactors[1320] = 00.000902;
scaleFactors[1319] = 00.000914;
scaleFactors[1318] = 00.000926;
scaleFactors[1317] = 00.000938;
scaleFactors[1316] = 00.000950;
scaleFactors[1315] = 00.000963;
scaleFactors[1314] = 00.000975;
scaleFactors[1313] = 00.000988;
scaleFactors[1312] = 00.001001;
scaleFactors[1311] = 00.001014;
scaleFactors[1310] = 00.001027;
scaleFactors[1309] = 00.001041;
scaleFactors[1308] = 00.001055;
scaleFactors[1307] = 00.001068;
scaleFactors[1306] = 00.001082;
scaleFactors[1305] = 00.001097;
scaleFactors[1304] = 00.001111;
scaleFactors[1303] = 00.001125;
scaleFactors[1302] = 00.001140;
scaleFactors[1301] = 00.001155;
scaleFactors[1300] = 00.001170;
scaleFactors[1299] = 00.001186;
scaleFactors[1298] = 00.001201;
scaleFactors[1297] = 00.001217;
scaleFactors[1296] = 00.001233;
scaleFactors[1295] = 00.001249;
scaleFactors[1294] = 00.001265;
scaleFactors[1293] = 00.001282;
scaleFactors[1292] = 00.001299;
scaleFactors[1291] = 00.001316;
scaleFactors[1290] = 00.001333;
scaleFactors[1289] = 00.001350;
scaleFactors[1288] = 00.001368;
scaleFactors[1287] = 00.001386;
scaleFactors[1286] = 00.001404;
scaleFactors[1285] = 00.001423;
scaleFactors[1284] = 00.001441;
scaleFactors[1283] = 00.001460;
scaleFactors[1282] = 00.001479;
scaleFactors[1281] = 00.001499;
scaleFactors[1280] = 00.001518;
scaleFactors[1279] = 00.001538;
scaleFactors[1278] = 00.001558;
scaleFactors[1277] = 00.001579;
scaleFactors[1276] = 00.001599;
scaleFactors[1275] = 00.001620;
scaleFactors[1274] = 00.001642;
scaleFactors[1273] = 00.001663;
scaleFactors[1272] = 00.001685;
scaleFactors[1271] = 00.001707;
scaleFactors[1270] = 00.001729;
scaleFactors[1269] = 00.001752;
scaleFactors[1268] = 00.001775;
scaleFactors[1267] = 00.001798;
scaleFactors[1266] = 00.001822;
scaleFactors[1265] = 00.001846;
scaleFactors[1264] = 00.001870;
scaleFactors[1263] = 00.001894;
scaleFactors[1262] = 00.001919;
scaleFactors[1261] = 00.001944;
scaleFactors[1260] = 00.001970;
scaleFactors[1259] = 00.001995;
scaleFactors[1258] = 00.002022;
scaleFactors[1257] = 00.002048;
scaleFactors[1256] = 00.002075;
scaleFactors[1255] = 00.002102;
scaleFactors[1254] = 00.002130;
scaleFactors[1253] = 00.002157;
scaleFactors[1252] = 00.002186;
scaleFactors[1251] = 00.002214;
scaleFactors[1250] = 00.002243;
scaleFactors[1249] = 00.002273;
scaleFactors[1248] = 00.002303;
scaleFactors[1247] = 00.002333;
scaleFactors[1246] = 00.002363;
scaleFactors[1245] = 00.002394;
scaleFactors[1244] = 00.002426;
scaleFactors[1243] = 00.002457;
scaleFactors[1242] = 00.002490;
scaleFactors[1241] = 00.002522;
scaleFactors[1240] = 00.002555;
scaleFactors[1239] = 00.002589;
scaleFactors[1238] = 00.002623;
scaleFactors[1237] = 00.002657;
scaleFactors[1236] = 00.002692;
scaleFactors[1235] = 00.002727;
scaleFactors[1234] = 00.002763;
scaleFactors[1233] = 00.002799;
scaleFactors[1232] = 00.002836;
scaleFactors[1231] = 00.002873;
scaleFactors[1230] = 00.002910;
scaleFactors[1229] = 00.002949;
scaleFactors[1228] = 00.002987;
scaleFactors[1227] = 00.003026;
scaleFactors[1226] = 00.003066;
scaleFactors[1225] = 00.003106;
scaleFactors[1224] = 00.003147;
scaleFactors[1223] = 00.003188;
scaleFactors[1222] = 00.003230;
scaleFactors[1221] = 00.003272;
scaleFactors[1220] = 00.003315;
scaleFactors[1219] = 00.003358;
scaleFactors[1218] = 00.003402;
scaleFactors[1217] = 00.003447;
scaleFactors[1216] = 00.003492;
scaleFactors[1215] = 00.003538;
scaleFactors[1214] = 00.003584;
scaleFactors[1213] = 00.003631;
scaleFactors[1212] = 00.003679;
scaleFactors[1211] = 00.003727;
scaleFactors[1210] = 00.003776;
scaleFactors[1209] = 00.003825;
scaleFactors[1208] = 00.003875;
scaleFactors[1207] = 00.003926;
scaleFactors[1206] = 00.003977;
scaleFactors[1205] = 00.004030;
scaleFactors[1204] = 00.004082;
scaleFactors[1203] = 00.004136;
scaleFactors[1202] = 00.004190;
scaleFactors[1201] = 00.004245;
scaleFactors[1200] = 00.004301;
scaleFactors[1199] = 00.004357;
scaleFactors[1198] = 00.004414;
scaleFactors[1197] = 00.004472;
scaleFactors[1196] = 00.004530;
scaleFactors[1195] = 00.004590;
scaleFactors[1194] = 00.004650;
scaleFactors[1193] = 00.004711;
scaleFactors[1192] = 00.004772;
scaleFactors[1191] = 00.004835;
scaleFactors[1190] = 00.004898;
scaleFactors[1189] = 00.004962;
scaleFactors[1188] = 00.005027;
scaleFactors[1187] = 00.005093;
scaleFactors[1186] = 00.005160;
scaleFactors[1185] = 00.005228;
scaleFactors[1184] = 00.005296;
scaleFactors[1183] = 00.005366;
scaleFactors[1182] = 00.005436;
scaleFactors[1181] = 00.005507;
scaleFactors[1180] = 00.005579;
scaleFactors[1179] = 00.005652;
scaleFactors[1178] = 00.005726;
scaleFactors[1177] = 00.005801;
scaleFactors[1176] = 00.005877;
scaleFactors[1175] = 00.005954;
scaleFactors[1174] = 00.006032;
scaleFactors[1173] = 00.006111;
scaleFactors[1172] = 00.006191;
scaleFactors[1171] = 00.006272;
scaleFactors[1170] = 00.006355;
scaleFactors[1169] = 00.006438;
scaleFactors[1168] = 00.006522;
scaleFactors[1167] = 00.006608;
scaleFactors[1166] = 00.006694;
scaleFactors[1165] = 00.006782;
scaleFactors[1164] = 00.006871;
scaleFactors[1163] = 00.006961;
scaleFactors[1162] = 00.007052;
scaleFactors[1161] = 00.007144;
scaleFactors[1160] = 00.007238;
scaleFactors[1159] = 00.007333;
scaleFactors[1158] = 00.007429;
scaleFactors[1157] = 00.007526;
scaleFactors[1156] = 00.007625;
scaleFactors[1155] = 00.007725;
scaleFactors[1154] = 00.007826;
scaleFactors[1153] = 00.007928;
scaleFactors[1152] = 00.008032;
scaleFactors[1151] = 00.008137;
scaleFactors[1150] = 00.008244;
scaleFactors[1149] = 00.008352;
scaleFactors[1148] = 00.008461;
scaleFactors[1147] = 00.008572;
scaleFactors[1146] = 00.008685;
scaleFactors[1145] = 00.008798;
scaleFactors[1144] = 00.008914;
scaleFactors[1143] = 00.009030;
scaleFactors[1142] = 00.009149;
scaleFactors[1141] = 00.009269;
scaleFactors[1140] = 00.009390;
scaleFactors[1139] = 00.009513;
scaleFactors[1138] = 00.009638;
scaleFactors[1137] = 00.009764;
scaleFactors[1136] = 00.009892;
scaleFactors[1135] = 00.010021;
scaleFactors[1134] = 00.010153;
scaleFactors[1133] = 00.010286;
scaleFactors[1132] = 00.010420;
scaleFactors[1131] = 00.010557;
scaleFactors[1130] = 00.010695;
scaleFactors[1129] = 00.010835;
scaleFactors[1128] = 00.010977;
scaleFactors[1127] = 00.011121;
scaleFactors[1126] = 00.011267;
scaleFactors[1125] = 00.011414;
scaleFactors[1124] = 00.011564;
scaleFactors[1123] = 00.011715;
scaleFactors[1122] = 00.011869;
scaleFactors[1121] = 00.012024;
scaleFactors[1120] = 00.012182;
scaleFactors[1119] = 00.012341;
scaleFactors[1118] = 00.012503;
scaleFactors[1117] = 00.012667;
scaleFactors[1116] = 00.012833;
scaleFactors[1115] = 00.013001;
scaleFactors[1114] = 00.013171;
scaleFactors[1113] = 00.013344;
scaleFactors[1112] = 00.013518;
scaleFactors[1111] = 00.013696;
scaleFactors[1110] = 00.013875;
scaleFactors[1109] = 00.014057;
scaleFactors[1108] = 00.014241;
scaleFactors[1107] = 00.014427;
scaleFactors[1106] = 00.014616;
scaleFactors[1105] = 00.014808;
scaleFactors[1104] = 00.015002;
scaleFactors[1103] = 00.015198;
scaleFactors[1102] = 00.015398;
scaleFactors[1101] = 00.015599;
scaleFactors[1100] = 00.015804;
scaleFactors[1099] = 00.016011;
scaleFactors[1098] = 00.016220;
scaleFactors[1097] = 00.016433;
scaleFactors[1096] = 00.016648;
scaleFactors[1095] = 00.016866;
scaleFactors[1094] = 00.017087;
scaleFactors[1093] = 00.017311;
scaleFactors[1092] = 00.017538;
scaleFactors[1091] = 00.017767;
scaleFactors[1090] = 00.018000;
scaleFactors[1089] = 00.018236;
scaleFactors[1088] = 00.018475;
scaleFactors[1087] = 00.018717;
scaleFactors[1086] = 00.018962;
scaleFactors[1085] = 00.019211;
scaleFactors[1084] = 00.019462;
scaleFactors[1083] = 00.019717;
scaleFactors[1082] = 00.019975;
scaleFactors[1081] = 00.020237;
scaleFactors[1080] = 00.020502;
scaleFactors[1079] = 00.020771;
scaleFactors[1078] = 00.021043;
scaleFactors[1077] = 00.021319;
scaleFactors[1076] = 00.021598;
scaleFactors[1075] = 00.021881;
scaleFactors[1074] = 00.022167;
scaleFactors[1073] = 00.022458;
scaleFactors[1072] = 00.022752;
scaleFactors[1071] = 00.023050;
scaleFactors[1070] = 00.023352;
scaleFactors[1069] = 00.023658;
scaleFactors[1068] = 00.023968;
scaleFactors[1067] = 00.024282;
scaleFactors[1066] = 00.024600;
scaleFactors[1065] = 00.024922;
scaleFactors[1064] = 00.025249;
scaleFactors[1063] = 00.025579;
scaleFactors[1062] = 00.025915;
scaleFactors[1061] = 00.026254;
scaleFactors[1060] = 00.026598;
scaleFactors[1059] = 00.026946;
scaleFactors[1058] = 00.027299;
scaleFactors[1057] = 00.027657;
scaleFactors[1056] = 00.028019;
scaleFactors[1055] = 00.028386;
scaleFactors[1054] = 00.028758;
scaleFactors[1053] = 00.029135;
scaleFactors[1052] = 00.029517;
scaleFactors[1051] = 00.029903;
scaleFactors[1050] = 00.030295;
scaleFactors[1049] = 00.030692;
scaleFactors[1048] = 00.031094;
scaleFactors[1047] = 00.031501;
scaleFactors[1046] = 00.031914;
scaleFactors[1045] = 00.032332;
scaleFactors[1044] = 00.032756;
scaleFactors[1043] = 00.033185;
scaleFactors[1042] = 00.033619;
scaleFactors[1041] = 00.034060;
scaleFactors[1040] = 00.034506;
scaleFactors[1039] = 00.034958;
scaleFactors[1038] = 00.035416;
scaleFactors[1037] = 00.035880;
scaleFactors[1036] = 00.036350;
scaleFactors[1035] = 00.036826;
scaleFactors[1034] = 00.037309;
scaleFactors[1033] = 00.037797;
scaleFactors[1032] = 00.038292;
scaleFactors[1031] = 00.038794;
scaleFactors[1030] = 00.039302;
scaleFactors[1029] = 00.039817;
scaleFactors[1028] = 00.040339;
scaleFactors[1027] = 00.040867;
scaleFactors[1026] = 00.041403;
scaleFactors[1025] = 00.041945;
scaleFactors[1024] = 00.042494;
scaleFactors[1023] = 00.043051;
scaleFactors[1022] = 00.043615;
scaleFactors[1021] = 00.044186;
scaleFactors[1020] = 00.044765;
scaleFactors[1019] = 00.045352;
scaleFactors[1018] = 00.045946;
scaleFactors[1017] = 00.046548;
scaleFactors[1016] = 00.047157;
scaleFactors[1015] = 00.047775;
scaleFactors[1014] = 00.048401;
scaleFactors[1013] = 00.049035;
scaleFactors[1012] = 00.049677;
scaleFactors[1011] = 00.050328;
scaleFactors[1010] = 00.050988;
scaleFactors[1009] = 00.051656;
scaleFactors[1008] = 00.052332;
scaleFactors[1007] = 00.053018;
scaleFactors[1006] = 00.053712;
scaleFactors[1005] = 00.054416;
scaleFactors[1004] = 00.055129;
scaleFactors[1003] = 00.055851;
scaleFactors[1002] = 00.056583;
scaleFactors[1001] = 00.057324;
scaleFactors[1000] = 00.058075;
scaleFactors[999] = 00.058836;
scaleFactors[998] = 00.059606;
scaleFactors[997] = 00.060387;
scaleFactors[996] = 00.061178;
scaleFactors[995] = 00.061980;
scaleFactors[994] = 00.062792;
scaleFactors[993] = 00.063614;
scaleFactors[992] = 00.064448;
scaleFactors[991] = 00.065292;
scaleFactors[990] = 00.066147;
scaleFactors[989] = 00.067014;
scaleFactors[988] = 00.067892;
scaleFactors[987] = 00.068781;
scaleFactors[986] = 00.069682;
scaleFactors[985] = 00.070595;
scaleFactors[984] = 00.071520;
scaleFactors[983] = 00.072456;
scaleFactors[982] = 00.073406;
scaleFactors[981] = 00.074367;
scaleFactors[980] = 00.075342;
scaleFactors[979] = 00.076328;
scaleFactors[978] = 00.077328;
scaleFactors[977] = 00.078341;
scaleFactors[976] = 00.079368;
scaleFactors[975] = 00.080407;
scaleFactors[974] = 00.081461;
scaleFactors[973] = 00.082528;
scaleFactors[972] = 00.083609;
scaleFactors[971] = 00.084704;
scaleFactors[970] = 00.085814;
scaleFactors[969] = 00.086938;
scaleFactors[968] = 00.088077;
scaleFactors[967] = 00.089231;
scaleFactors[966] = 00.090400;
scaleFactors[965] = 00.091584;
scaleFactors[964] = 00.092784;
scaleFactors[963] = 00.093999;
scaleFactors[962] = 00.095231;
scaleFactors[961] = 00.096478;
scaleFactors[960] = 00.097742;
scaleFactors[959] = 00.099022;
scaleFactors[958] = 00.100320;
scaleFactors[957] = 00.101634;
scaleFactors[956] = 00.102965;
scaleFactors[955] = 00.104314;
scaleFactors[954] = 00.105680;
scaleFactors[953] = 00.107065;
scaleFactors[952] = 00.108467;
scaleFactors[951] = 00.109888;
scaleFactors[950] = 00.111328;
scaleFactors[949] = 00.112786;
scaleFactors[948] = 00.114264;
scaleFactors[947] = 00.115761;
scaleFactors[946] = 00.117277;
scaleFactors[945] = 00.118813;
scaleFactors[944] = 00.120370;
scaleFactors[943] = 00.121947;
scaleFactors[942] = 00.123544;
scaleFactors[941] = 00.125163;
scaleFactors[940] = 00.126802;
scaleFactors[939] = 00.128464;
scaleFactors[938] = 00.130146;
scaleFactors[937] = 00.131851;
scaleFactors[936] = 00.133579;
scaleFactors[935] = 00.135328;
scaleFactors[934] = 00.137101;
scaleFactors[933] = 00.138897;
scaleFactors[932] = 00.140717;
scaleFactors[931] = 00.142560;
scaleFactors[930] = 00.144428;
scaleFactors[929] = 00.146320;
scaleFactors[928] = 00.148237;
scaleFactors[927] = 00.150178;
scaleFactors[926] = 00.152146;
scaleFactors[925] = 00.154139;
scaleFactors[924] = 00.156158;
scaleFactors[923] = 00.158204;
scaleFactors[922] = 00.160276;
scaleFactors[921] = 00.162376;
scaleFactors[920] = 00.164503;
scaleFactors[919] = 00.166658;
scaleFactors[918] = 00.168841;
scaleFactors[917] = 00.171053;
scaleFactors[916] = 00.173294;
scaleFactors[915] = 00.175564;
scaleFactors[914] = 00.177864;
scaleFactors[913] = 00.180194;
scaleFactors[912] = 00.182555;
scaleFactors[911] = 00.184946;
scaleFactors[910] = 00.187369;
scaleFactors[909] = 00.189823;
scaleFactors[908] = 00.192310;
scaleFactors[907] = 00.194829;
scaleFactors[906] = 00.197382;
scaleFactors[905] = 00.199967;
scaleFactors[904] = 00.202587;
scaleFactors[903] = 00.205241;
scaleFactors[902] = 00.207929;
scaleFactors[901] = 00.210653;
scaleFactors[900] = 00.213413;
scaleFactors[899] = 00.216209;
scaleFactors[898] = 00.219041;
scaleFactors[897] = 00.221910;
scaleFactors[896] = 00.224817;
scaleFactors[895] = 00.227763;
scaleFactors[894] = 00.230746;
scaleFactors[893] = 00.233769;
scaleFactors[892] = 00.236831;
scaleFactors[891] = 00.239934;
scaleFactors[890] = 00.243077;
scaleFactors[889] = 00.246261;
scaleFactors[888] = 00.249487;
scaleFactors[887] = 00.252756;
scaleFactors[886] = 00.256067;
scaleFactors[885] = 00.259421;
scaleFactors[884] = 00.262820;
scaleFactors[883] = 00.266263;
scaleFactors[882] = 00.269751;
scaleFactors[881] = 00.273284;
scaleFactors[880] = 00.276864;
scaleFactors[879] = 00.280491;
scaleFactors[878] = 00.284166;
scaleFactors[877] = 00.287888;
scaleFactors[876] = 00.291660;
scaleFactors[875] = 00.295480;
scaleFactors[874] = 00.299351;
scaleFactors[873] = 00.303273;
scaleFactors[872] = 00.307246;
scaleFactors[871] = 00.311271;
scaleFactors[870] = 00.315348;
scaleFactors[869] = 00.319479;
scaleFactors[868] = 00.323665;
scaleFactors[867] = 00.327905;
scaleFactors[866] = 00.332200;
scaleFactors[865] = 00.336552;
scaleFactors[864] = 00.340961;
scaleFactors[863] = 00.345427;
scaleFactors[862] = 00.349952;
scaleFactors[861] = 00.354537;
scaleFactors[860] = 00.359181;
scaleFactors[859] = 00.363887;
scaleFactors[858] = 00.368653;
scaleFactors[857] = 00.373483;
scaleFactors[856] = 00.378375;
scaleFactors[855] = 00.383332;
scaleFactors[854] = 00.388354;
scaleFactors[853] = 00.393441;
scaleFactors[852] = 00.398595;
scaleFactors[851] = 00.403817;
scaleFactors[850] = 00.409107;
scaleFactors[849] = 00.414466;
scaleFactors[848] = 00.419896;
scaleFactors[847] = 00.425396;
scaleFactors[846] = 00.430969;
scaleFactors[845] = 00.436615;
scaleFactors[844] = 00.442335;
scaleFactors[843] = 00.448129;
scaleFactors[842] = 00.454000;
scaleFactors[841] = 00.459947;
scaleFactors[840] = 00.465972;
scaleFactors[839] = 00.472077;
scaleFactors[838] = 00.478261;
scaleFactors[837] = 00.484526;
scaleFactors[836] = 00.490873;
scaleFactors[835] = 00.497304;
scaleFactors[834] = 00.503819;
scaleFactors[833] = 00.510419;
scaleFactors[832] = 00.517105;
scaleFactors[831] = 00.523879;
scaleFactors[830] = 00.530742;
scaleFactors[829] = 00.537695;
scaleFactors[828] = 00.544739;
scaleFactors[827] = 00.551875;
scaleFactors[826] = 00.559104;
scaleFactors[825] = 00.566428;
scaleFactors[824] = 00.573849;
scaleFactors[823] = 00.581366;
scaleFactors[822] = 00.588982;
scaleFactors[821] = 00.596698;
scaleFactors[820] = 00.604515;
scaleFactors[819] = 00.612434;
scaleFactors[818] = 00.620457;
scaleFactors[817] = 00.628585;
scaleFactors[816] = 00.636819;
scaleFactors[815] = 00.645161;
scaleFactors[814] = 00.653613;
scaleFactors[813] = 00.662175;
scaleFactors[812] = 00.670850;
scaleFactors[811] = 00.679638;
scaleFactors[810] = 00.688541;
scaleFactors[809] = 00.697561;
scaleFactors[808] = 00.706699;
scaleFactors[807] = 00.715957;
scaleFactors[806] = 00.725336;
scaleFactors[805] = 00.734838;
scaleFactors[804] = 00.744464;
scaleFactors[803] = 00.754217;
scaleFactors[802] = 00.764097;
scaleFactors[801] = 00.774107;
scaleFactors[800] = 00.784248;
scaleFactors[799] = 00.794521;
scaleFactors[798] = 00.804930;
scaleFactors[797] = 00.815474;
scaleFactors[796] = 00.826157;
scaleFactors[795] = 00.836980;
scaleFactors[794] = 00.847944;
scaleFactors[793] = 00.859052;
scaleFactors[792] = 00.870306;
scaleFactors[791] = 00.881707;
scaleFactors[790] = 00.893257;
scaleFactors[789] = 00.904959;
scaleFactors[788] = 00.916814;
scaleFactors[787] = 00.928824;
scaleFactors[786] = 00.940992;
scaleFactors[785] = 00.953319;
scaleFactors[784] = 00.965807;
scaleFactors[783] = 00.978459;
scaleFactors[782] = 00.991277;
scaleFactors[781] = 1.004263;
scaleFactors[780] = 1.017419;
scaleFactors[779] = 1.030747;
scaleFactors[778] = 1.044250;
scaleFactors[777] = 1.057930;
scaleFactors[776] = 1.071789;
scaleFactors[775] = 1.085829;
scaleFactors[774] = 1.100053;
scaleFactors[773] = 1.114464;
scaleFactors[772] = 1.129064;
scaleFactors[771] = 1.143854;
scaleFactors[770] = 1.158839;
scaleFactors[769] = 1.174020;
scaleFactors[768] = 1.189399;
scaleFactors[767] = 1.204981;
scaleFactors[766] = 1.220766;
scaleFactors[765] = 1.236758;
scaleFactors[764] = 1.252960;
scaleFactors[763] = 1.269373;
scaleFactors[762] = 1.286002;
scaleFactors[761] = 1.302849;
scaleFactors[760] = 1.319916;
scaleFactors[759] = 1.337207;
scaleFactors[758] = 1.354725;
scaleFactors[757] = 1.372472;
scaleFactors[756] = 1.390451;
scaleFactors[755] = 1.408666;
scaleFactors[754] = 1.427119;
scaleFactors[753] = 1.445815;
scaleFactors[752] = 1.464755;
scaleFactors[751] = 1.483943;
scaleFactors[750] = 1.503383;
scaleFactors[749] = 1.523077;
scaleFactors[748] = 1.543030;
scaleFactors[747] = 1.563243;
scaleFactors[746] = 1.583722;
scaleFactors[745] = 1.604469;
scaleFactors[744] = 1.625487;
scaleFactors[743] = 1.646781;
scaleFactors[742] = 1.668354;
scaleFactors[741] = 1.690210;
scaleFactors[740] = 1.712351;
scaleFactors[739] = 1.734783;
scaleFactors[738] = 1.757509;
scaleFactors[737] = 1.780532;
scaleFactors[736] = 1.803857;
scaleFactors[735] = 1.827488;
scaleFactors[734] = 1.851428;
scaleFactors[733] = 1.875682;
scaleFactors[732] = 1.900253;
scaleFactors[731] = 1.925147;
scaleFactors[730] = 1.950366;
scaleFactors[729] = 1.975916;
scaleFactors[728] = 2.001801;
scaleFactors[727] = 2.028024;
scaleFactors[726] = 2.054591;
scaleFactors[725] = 2.081507;
scaleFactors[724] = 2.108774;
scaleFactors[723] = 2.136400;
scaleFactors[722] = 2.164387;
scaleFactors[721] = 2.192740;
scaleFactors[720] = 2.221465;
scaleFactors[719] = 2.250566;
scaleFactors[718] = 2.280048;
scaleFactors[717] = 2.309917;
scaleFactors[716] = 2.340177;
scaleFactors[715] = 2.370833;
scaleFactors[714] = 2.401891;
scaleFactors[713] = 2.433356;
scaleFactors[712] = 2.465233;
scaleFactors[711] = 2.497528;
scaleFactors[710] = 2.530246;
scaleFactors[709] = 2.563392;
scaleFactors[708] = 2.596972;
scaleFactors[707] = 2.630993;
scaleFactors[706] = 2.665459;
scaleFactors[705] = 2.700377;
scaleFactors[704] = 2.735752;
scaleFactors[703] = 2.771590;
scaleFactors[702] = 2.807898;
scaleFactors[701] = 2.844681;
scaleFactors[700] = 2.881947;
scaleFactors[699] = 2.919700;
scaleFactors[698] = 2.957948;
scaleFactors[697] = 2.996697;
scaleFactors[696] = 3.035954;
scaleFactors[695] = 3.075725;
scaleFactors[694] = 3.116017;
scaleFactors[693] = 3.156837;
scaleFactors[692] = 3.198192;
scaleFactors[691] = 3.240088;
scaleFactors[690] = 3.282533;
scaleFactors[689] = 3.325535;
scaleFactors[688] = 3.369099;
scaleFactors[687] = 3.413234;
scaleFactors[686] = 3.457948;
scaleFactors[685] = 3.503247;
scaleFactors[684] = 3.549140;
scaleFactors[683] = 3.595634;
scaleFactors[682] = 3.642737;
scaleFactors[681] = 3.690457;
scaleFactors[680] = 3.738802;
scaleFactors[679] = 3.787780;
scaleFactors[678] = 3.837400;
scaleFactors[677] = 3.887670;
scaleFactors[676] = 3.938599;
scaleFactors[675] = 3.990194;
scaleFactors[674] = 4.042466;
scaleFactors[673] = 4.095423;
scaleFactors[672] = 4.149073;
scaleFactors[671] = 4.203426;
scaleFactors[670] = 4.258491;
scaleFactors[669] = 4.314277;
scaleFactors[668] = 4.370794;
scaleFactors[667] = 4.428052;
scaleFactors[666] = 4.486060;
scaleFactors[665] = 4.544827;
scaleFactors[664] = 4.604364;
scaleFactors[663] = 4.664682;
scaleFactors[662] = 4.725790;
scaleFactors[661] = 4.787697;
scaleFactors[660] = 4.850416;
scaleFactors[659] = 4.913957;
scaleFactors[658] = 4.978330;
scaleFactors[657] = 5.043546;
scaleFactors[656] = 5.109616;
scaleFactors[655] = 5.176552;
scaleFactors[654] = 5.244365;
scaleFactors[653] = 5.313066;
scaleFactors[652] = 5.382668;
scaleFactors[651] = 5.453181;
scaleFactors[650] = 5.524618;
scaleFactors[649] = 5.596991;
scaleFactors[648] = 5.670311;
scaleFactors[647] = 5.744593;
scaleFactors[646] = 5.819847;
scaleFactors[645] = 5.896087;
scaleFactors[644] = 5.973326;
scaleFactors[643] = 6.051577;
scaleFactors[642] = 6.130853;
scaleFactors[641] = 6.211167;
scaleFactors[640] = 6.292533;
scaleFactors[639] = 6.374966;
scaleFactors[638] = 6.458478;
scaleFactors[637] = 6.543084;
scaleFactors[636] = 6.628799;
scaleFactors[635] = 6.715636;
scaleFactors[634] = 6.803611;
scaleFactors[633] = 6.892739;
scaleFactors[632] = 6.983034;
scaleFactors[631] = 7.074512;
scaleFactors[630] = 7.167188;
scaleFactors[629] = 7.261078;
scaleFactors[628] = 7.356198;
scaleFactors[627] = 7.452565;
scaleFactors[626] = 7.550193;
scaleFactors[625] = 7.649101;
scaleFactors[624] = 7.749305;
scaleFactors[623] = 7.850821;
scaleFactors[622] = 7.953667;
scaleFactors[621] = 8.057860;
scaleFactors[620] = 8.163419;
scaleFactors[619] = 8.270360;
scaleFactors[618] = 8.378702;
scaleFactors[617] = 8.488463;
scaleFactors[616] = 8.599663;
scaleFactors[615] = 8.712318;
scaleFactors[614] = 8.826450;
scaleFactors[613] = 8.942077;
scaleFactors[612] = 9.059218;
scaleFactors[611] = 9.177895;
scaleFactors[610] = 9.298125;
scaleFactors[609] = 9.419931;
scaleFactors[608] = 9.543333;
scaleFactors[607] = 9.668351;
scaleFactors[606] = 9.795007;
scaleFactors[605] = 9.923322;
scaleFactors[604] = 10.053317;
scaleFactors[603] = 10.185016;
scaleFactors[602] = 10.318439;
scaleFactors[601] = 10.453611;
scaleFactors[600] = 10.590554;
scaleFactors[599] = 10.729291;
scaleFactors[598] = 10.869845;
scaleFactors[597] = 11.012240;
scaleFactors[596] = 11.156501;
scaleFactors[595] = 11.302651;
scaleFactors[594] = 11.450716;
scaleFactors[593] = 11.600720;
scaleFactors[592] = 11.752690;
scaleFactors[591] = 11.906651;
scaleFactors[590] = 12.062628;
scaleFactors[589] = 12.220649;
scaleFactors[588] = 12.380739;
scaleFactors[587] = 12.542927;
scaleFactors[586] = 12.707239;
scaleFactors[585] = 12.873704;
scaleFactors[584] = 13.042350;
scaleFactors[583] = 13.213205;
scaleFactors[582] = 13.386299;
scaleFactors[581] = 13.561660;
scaleFactors[580] = 13.739318;
scaleFactors[579] = 13.919303;
scaleFactors[578] = 14.101646;
scaleFactors[577] = 14.286379;
scaleFactors[576] = 14.473531;
scaleFactors[575] = 14.663135;
scaleFactors[574] = 14.855222;
scaleFactors[573] = 15.049826;
scaleFactors[572] = 15.246979;
scaleFactors[571] = 15.446714;
scaleFactors[570] = 15.649067;
scaleFactors[569] = 15.854070;
scaleFactors[568] = 16.061758;
scaleFactors[567] = 16.272167;
scaleFactors[566] = 16.485332;
scaleFactors[565] = 16.701290;
scaleFactors[564] = 16.920078;
scaleFactors[563] = 17.141731;
scaleFactors[562] = 17.366289;
scaleFactors[561] = 17.593788;
scaleFactors[560] = 17.824266;
scaleFactors[559] = 18.057764;
scaleFactors[558] = 18.294321;
scaleFactors[557] = 18.533978;
scaleFactors[556] = 18.776773;
scaleFactors[555] = 19.022749;
scaleFactors[554] = 19.271948;
scaleFactors[553] = 19.524410;
scaleFactors[552] = 19.780180;
scaleFactors[551] = 20.039301;
scaleFactors[550] = 20.301817;
scaleFactors[549] = 20.567772;
scaleFactors[548] = 20.837210;
scaleFactors[547] = 21.110178;
scaleFactors[546] = 21.386723;
scaleFactors[545] = 21.666889;
scaleFactors[544] = 21.950726;
scaleFactors[543] = 22.238281;
scaleFactors[542] = 22.529604;
scaleFactors[541] = 22.824743;
scaleFactors[540] = 23.123749;
scaleFactors[539] = 23.426670;
scaleFactors[538] = 23.733561;
scaleFactors[537] = 24.044472;
scaleFactors[536] = 24.359455;
scaleFactors[535] = 24.678564;
scaleFactors[534] = 25.001854;
scaleFactors[533] = 25.329378;
scaleFactors[532] = 25.661194;
scaleFactors[531] = 25.997356;
scaleFactors[530] = 26.337923;
scaleFactors[529] = 26.682951;
scaleFactors[528] = 27.032499;
scaleFactors[527] = 27.386625;
scaleFactors[526] = 27.745390;
scaleFactors[525] = 28.108856;
scaleFactors[524] = 28.477083;
scaleFactors[523] = 28.850134;
scaleFactors[522] = 29.228071;
scaleFactors[521] = 29.610960;
scaleFactors[520] = 29.998865;
scaleFactors[519] = 30.391851;
scaleFactors[518] = 30.789986;
scaleFactors[517] = 31.193335;
scaleFactors[516] = 31.601969;
scaleFactors[515] = 32.015957;
scaleFactors[514] = 32.435368;
scaleFactors[513] = 32.860271;
scaleFactors[512] = 33.290741;
scaleFactors[511] = 33.726852;
scaleFactors[510] = 34.168674;
scaleFactors[509] = 34.616283;
scaleFactors[508] = 35.069759;
scaleFactors[507] = 35.529175;
scaleFactors[506] = 35.994610;
scaleFactors[505] = 36.466141;
scaleFactors[504] = 36.943848;
scaleFactors[503] = 37.427814;
scaleFactors[502] = 37.918121;
scaleFactors[501] = 38.414848;
scaleFactors[500] = 38.918083;
scaleFactors[499] = 39.427910;
scaleFactors[498] = 39.944416;
scaleFactors[497] = 40.467690;
scaleFactors[496] = 40.997818;
scaleFactors[495] = 41.534889;
scaleFactors[494] = 42.078999;
scaleFactors[493] = 42.630234;
scaleFactors[492] = 43.188690;
scaleFactors[491] = 43.754463;
scaleFactors[490] = 44.327648;
scaleFactors[489] = 44.908340;
scaleFactors[488] = 45.496639;
scaleFactors[487] = 46.092648;
scaleFactors[486] = 46.696461;
scaleFactors[485] = 47.308186;
scaleFactors[484] = 47.927925;
scaleFactors[483] = 48.555782;
scaleFactors[482] = 49.191864;
scaleFactors[481] = 49.836277;
scaleFactors[480] = 50.489132;
scaleFactors[479] = 51.150539;
scaleFactors[478] = 51.820614;
scaleFactors[477] = 52.499466;
scaleFactors[476] = 53.187210;
scaleFactors[475] = 53.883965;
scaleFactors[474] = 54.589848;
scaleFactors[473] = 55.304977;
scaleFactors[472] = 56.029472;
scaleFactors[471] = 56.763458;
scaleFactors[470] = 57.507061;
scaleFactors[469] = 58.260406;
scaleFactors[468] = 59.023621;
scaleFactors[467] = 59.796833;
scaleFactors[466] = 60.580173;
scaleFactors[465] = 61.373775;
scaleFactors[464] = 62.177773;
scaleFactors[463] = 62.992302;
scaleFactors[462] = 63.817501;
scaleFactors[461] = 64.653511;
scaleFactors[460] = 65.500473;
scaleFactors[459] = 66.358528;
scaleFactors[458] = 67.227829;
scaleFactors[457] = 68.108513;
scaleFactors[456] = 69.000740;
scaleFactors[455] = 69.904655;
scaleFactors[454] = 70.820412;
scaleFactors[453] = 71.748161;
scaleFactors[452] = 72.688065;
scaleFactors[451] = 73.640282;
scaleFactors[450] = 74.604973;
scaleFactors[449] = 75.582298;
scaleFactors[448] = 76.572426;
scaleFactors[447] = 77.575523;
scaleFactors[446] = 78.591766;
scaleFactors[445] = 79.621323;
scaleFactors[444] = 80.664368;
scaleFactors[443] = 81.721077;
scaleFactors[442] = 82.791626;
scaleFactors[441] = 83.876198;
scaleFactors[440] = 84.974976;
scaleFactors[439] = 86.088150;
scaleFactors[438] = 87.215904;
scaleFactors[437] = 88.358437;
scaleFactors[436] = 89.515938;
scaleFactors[435] = 90.688599;
scaleFactors[434] = 91.876625;
scaleFactors[433] = 93.080208;
scaleFactors[432] = 94.299561;
scaleFactors[431] = 95.534889;
scaleFactors[430] = 96.786400;
scaleFactors[429] = 98.054306;
scaleFactors[428] = 99.338821;
scaleFactors[427] = 100.640160;
scaleFactors[426] = 101.958549;
scaleFactors[425] = 103.294212;
scaleFactors[424] = 104.647369;
scaleFactors[423] = 106.018250;
scaleFactors[422] = 107.407089;
scaleFactors[421] = 108.814125;
scaleFactors[420] = 110.239594;
scaleFactors[419] = 111.683739;
scaleFactors[418] = 113.146797;
scaleFactors[417] = 114.629021;
scaleFactors[416] = 116.130661;
scaleFactors[415] = 117.651978;
scaleFactors[414] = 119.193222;
scaleFactors[413] = 120.754654;
scaleFactors[412] = 122.336540;
scaleFactors[411] = 123.939156;
scaleFactors[410] = 125.562759;
scaleFactors[409] = 127.207634;
scaleFactors[408] = 128.874054;
scaleFactors[407] = 130.562302;
scaleFactors[406] = 132.272675;
scaleFactors[405] = 134.005447;
scaleFactors[404] = 135.760925;
scaleFactors[403] = 137.539398;
scaleFactors[402] = 139.341171;
scaleFactors[401] = 141.166550;
scaleFactors[400] = 143.015839;
scaleFactors[399] = 144.889343;
scaleFactors[398] = 146.787399;
scaleFactors[397] = 148.710312;
scaleFactors[396] = 150.658417;
scaleFactors[395] = 152.632050;
scaleFactors[394] = 154.631531;
scaleFactors[393] = 156.657211;
scaleFactors[392] = 158.709427;
scaleFactors[391] = 160.788528;
scaleFactors[390] = 162.894867;
scaleFactors[389] = 165.028793;
scaleFactors[388] = 167.190674;
scaleFactors[387] = 169.380875;
scaleFactors[386] = 171.599762;
scaleFactors[385] = 173.847717;
scaleFactors[384] = 176.125122;
scaleFactors[383] = 178.432373;
scaleFactors[382] = 180.769836;
scaleFactors[381] = 183.137924;
scaleFactors[380] = 185.537033;
scaleFactors[379] = 187.967575;
scaleFactors[378] = 190.429962;
scaleFactors[377] = 192.924606;
scaleFactors[376] = 195.451920;
scaleFactors[375] = 198.012344;
scaleFactors[374] = 200.606308;
scaleFactors[373] = 203.234253;
scaleFactors[372] = 205.896622;
scaleFactors[371] = 208.593872;
scaleFactors[370] = 211.326462;
scaleFactors[369] = 214.094849;
scaleFactors[368] = 216.899490;
scaleFactors[367] = 219.740875;
scaleFactors[366] = 222.619492;
scaleFactors[365] = 225.535812;
scaleFactors[364] = 228.490341;
scaleFactors[363] = 231.483566;
scaleFactors[362] = 234.516006;
scaleFactors[361] = 237.588165;
scaleFactors[360] = 240.700577;
scaleFactors[359] = 243.853760;
scaleFactors[358] = 247.048248;
scaleFactors[357] = 250.284592;
scaleFactors[356] = 253.563324;
scaleFactors[355] = 256.885010;
scaleFactors[354] = 260.250214;
scaleFactors[353] = 263.659485;
scaleFactors[352] = 267.113434;
scaleFactors[351] = 270.612640;
scaleFactors[350] = 274.157684;
scaleFactors[349] = 277.749146;
scaleFactors[348] = 281.387665;
scaleFactors[347] = 285.073853;
scaleFactors[346] = 288.808319;
scaleFactors[345] = 292.591705;
scaleFactors[344] = 296.424652;
scaleFactors[343] = 300.307831;
scaleFactors[342] = 304.241882;
scaleFactors[341] = 308.227448;
scaleFactors[340] = 312.265228;
scaleFactors[339] = 316.355927;
scaleFactors[338] = 320.500183;
scaleFactors[337] = 324.698730;
scaleFactors[336] = 328.952301;
scaleFactors[335] = 333.261597;
scaleFactors[334] = 337.627319;
scaleFactors[333] = 342.050232;
scaleFactors[332] = 346.531097;
scaleFactors[331] = 351.070679;
scaleFactors[330] = 355.669708;
scaleFactors[329] = 360.328979;
scaleFactors[328] = 365.049286;
scaleFactors[327] = 369.831451;
scaleFactors[326] = 374.676239;
scaleFactors[325] = 379.584503;
scaleFactors[324] = 384.557068;
scaleFactors[323] = 389.594788;
scaleFactors[322] = 394.698486;
scaleFactors[321] = 399.869049;
scaleFactors[320] = 405.107330;
scaleFactors[319] = 410.414246;
scaleFactors[318] = 415.790680;
scaleFactors[317] = 421.237549;
scaleFactors[316] = 426.755768;
scaleFactors[315] = 432.346283;
scaleFactors[314] = 438.010040;
scaleFactors[313] = 443.747986;
scaleFactors[312] = 449.561096;
scaleFactors[311] = 455.450348;
scaleFactors[310] = 461.416748;
scaleFactors[309] = 467.461334;
scaleFactors[308] = 473.585083;
scaleFactors[307] = 479.789062;
scaleFactors[306] = 486.074310;
scaleFactors[305] = 492.441895;
scaleFactors[304] = 498.892883;
scaleFactors[303] = 505.428406;
scaleFactors[302] = 512.049561;
scaleFactors[301] = 518.757446;
scaleFactors[300] = 525.553162;
scaleFactors[299] = 532.437927;
scaleFactors[298] = 539.412903;
scaleFactors[297] = 546.479248;
scaleFactors[296] = 553.638123;
scaleFactors[295] = 560.890808;
scaleFactors[294] = 568.238464;
scaleFactors[293] = 575.682434;
scaleFactors[292] = 583.223877;
scaleFactors[291] = 590.864136;
scaleFactors[290] = 598.604492;
scaleFactors[289] = 606.446228;
scaleFactors[288] = 614.390686;
scaleFactors[287] = 622.439209;
scaleFactors[286] = 630.593201;
scaleFactors[285] = 638.854004;
scaleFactors[284] = 647.223022;
scaleFactors[283] = 655.701660;
scaleFactors[282] = 664.291382;
scaleFactors[281] = 672.993591;
scaleFactors[280] = 681.809814;
scaleFactors[279] = 690.741516;
scaleFactors[278] = 699.790222;
scaleFactors[277] = 708.957520;
scaleFactors[276] = 718.244873;
scaleFactors[275] = 727.653931;
scaleFactors[274] = 737.186218;
scaleFactors[273] = 746.843384;
scaleFactors[272] = 756.627075;
scaleFactors[271] = 766.538940;
scaleFactors[270] = 776.580627;
scaleFactors[269] = 786.753845;
scaleFactors[268] = 797.060364;
scaleFactors[267] = 807.501892;
scaleFactors[266] = 818.080200;
scaleFactors[265] = 828.797058;
scaleFactors[264] = 839.654297;
scaleFactors[263] = 850.653809;
scaleFactors[262] = 861.797424;
scaleFactors[261] = 873.086975;
scaleFactors[260] = 884.524414;
scaleFactors[259] = 896.111694;
scaleFactors[258] = 907.850769;
scaleFactors[257] = 919.743652;
scaleFactors[256] = 931.792297;
scaleFactors[255] = 943.998779;
scaleFactors[254] = 956.365173;
scaleFactors[253] = 968.893555;
scaleFactors[252] = 981.586060;
scaleFactors[251] = 994.444885;
scaleFactors[250] = 1007.472168;
scaleFactors[249] = 1020.670105;
scaleFactors[248] = 1034.040894;
scaleFactors[247] = 1000.0;
scaleFactors[246] = 1000.0;
scaleFactors[245] = 1000.0;
scaleFactors[244] = 1000.0;
scaleFactors[243] = 1000.0;
scaleFactors[242] = 1000.0;
scaleFactors[241] = 1000.0;
scaleFactors[240] = 1000.0;
scaleFactors[239] = 1000.0;
scaleFactors[238] = 1000.0;
scaleFactors[237] = 1000.0;
scaleFactors[236] = 1000.0;
scaleFactors[235] = 1000.0;
scaleFactors[234] = 1000.0;
scaleFactors[233] = 1000.0;
scaleFactors[232] = 1000.0;
scaleFactors[231] = 1000.0;
scaleFactors[230] = 1000.0;
scaleFactors[229] = 1000.0;
scaleFactors[228] = 1000.0;
scaleFactors[227] = 1000.0;
scaleFactors[226] = 1000.0;
scaleFactors[225] = 1000.0;
scaleFactors[224] = 1000.0;
scaleFactors[223] = 1000.0;
scaleFactors[222] = 1000.0;
scaleFactors[221] = 1000.0;
scaleFactors[220] = 1000.0;
scaleFactors[219] = 1000.0;
scaleFactors[218] = 1000.0;
scaleFactors[217] = 1000.0;
scaleFactors[216] = 1000.0;
scaleFactors[215] = 1000.0;
scaleFactors[214] = 1000.0;
scaleFactors[213] = 1000.0;
scaleFactors[212] = 1000.0;
scaleFactors[211] = 1000.0;
scaleFactors[210] = 1000.0;
scaleFactors[209] = 1000.0;
scaleFactors[208] = 1000.0;
scaleFactors[207] = 1000.0;
scaleFactors[206] = 1000.0;
scaleFactors[205] = 1000.0;
scaleFactors[204] = 1000.0;
scaleFactors[203] = 1000.0;
scaleFactors[202] = 1000.0;
scaleFactors[201] = 1000.0;
scaleFactors[200] = 1000.0;
scaleFactors[199] = 1000.0;
scaleFactors[198] = 1000.0;
scaleFactors[197] = 1000.0;
scaleFactors[196] = 1000.0;
scaleFactors[195] = 1000.0;
scaleFactors[194] = 1000.0;
scaleFactors[193] = 1000.0;
scaleFactors[192] = 1000.0;
scaleFactors[191] = 1000.0;
scaleFactors[190] = 1000.0;
scaleFactors[189] = 1000.0;
scaleFactors[188] = 1000.0;
scaleFactors[187] = 1000.0;
scaleFactors[186] = 1000.0;
scaleFactors[185] = 1000.0;
scaleFactors[184] = 1000.0;
scaleFactors[183] = 1000.0;
scaleFactors[182] = 1000.0;
scaleFactors[181] = 1000.0;
scaleFactors[180] = 1000.0;
scaleFactors[179] = 1000.0;
scaleFactors[178] = 1000.0;
scaleFactors[177] = 1000.0;
scaleFactors[176] = 1000.0;
scaleFactors[175] = 1000.0;
scaleFactors[174] = 1000.0;
scaleFactors[173] = 1000.0;
scaleFactors[172] = 1000.0;
scaleFactors[171] = 1000.0;
scaleFactors[170] = 1000.0;
scaleFactors[169] = 1000.0;
scaleFactors[168] = 1000.0;
scaleFactors[167] = 1000.0;
scaleFactors[166] = 1000.0;
scaleFactors[165] = 1000.0;
scaleFactors[164] = 1000.0;
scaleFactors[163] = 1000.0;
scaleFactors[162] = 1000.0;
scaleFactors[161] = 1000.0;
scaleFactors[160] = 1000.0;
scaleFactors[159] = 1000.0;
scaleFactors[158] = 1000.0;
scaleFactors[157] = 1000.0;
scaleFactors[156] = 1000.0;
scaleFactors[155] = 1000.0;
scaleFactors[154] = 1000.0;
scaleFactors[153] = 1000.0;
scaleFactors[152] = 1000.0;
scaleFactors[151] = 1000.0;
scaleFactors[150] = 1000.0;
scaleFactors[149] = 1000.0;
scaleFactors[148] = 1000.0;
scaleFactors[147] = 1000.0;
scaleFactors[146] = 1000.0;
scaleFactors[145] = 1000.0;
scaleFactors[144] = 1000.0;
scaleFactors[143] = 1000.0;
scaleFactors[142] = 1000.0;
scaleFactors[141] = 1000.0;
scaleFactors[140] = 1000.0;
scaleFactors[139] = 1000.0;
scaleFactors[138] = 1000.0;
scaleFactors[137] = 1000.0;
scaleFactors[136] = 1000.0;
scaleFactors[135] = 1000.0;
scaleFactors[134] = 1000.0;
scaleFactors[133] = 1000.0;
scaleFactors[132] = 1000.0;
scaleFactors[131] = 1000.0;
scaleFactors[130] = 1000.0;
scaleFactors[129] = 1000.0;
scaleFactors[128] = 1000.0;
scaleFactors[127] = 1000.0;
scaleFactors[126] = 1000.0;
scaleFactors[125] = 1000.0;
scaleFactors[124] = 1000.0;
scaleFactors[123] = 1000.0;
scaleFactors[122] = 1000.0;
scaleFactors[121] = 1000.0;
scaleFactors[120] = 1000.0;
scaleFactors[119] = 1000.0;
scaleFactors[118] = 1000.0;
scaleFactors[117] = 1000.0;
scaleFactors[116] = 1000.0;
scaleFactors[115] = 1000.0;
scaleFactors[114] = 1000.0;
scaleFactors[113] = 1000.0;
scaleFactors[112] = 1000.0;
scaleFactors[111] = 1000.0;
scaleFactors[110] = 1000.0;
scaleFactors[109] = 1000.0;
scaleFactors[108] = 1000.0;
scaleFactors[107] = 1000.0;
scaleFactors[106] = 1000.0;
scaleFactors[105] = 1000.0;
scaleFactors[104] = 1000.0;
scaleFactors[103] = 1000.0;
scaleFactors[102] = 1000.0;
scaleFactors[101] = 1000.0;
scaleFactors[100] = 1000.0;
scaleFactors[99] = 1000.0;
scaleFactors[98] = 1000.0;
scaleFactors[97] = 1000.0;
scaleFactors[96] = 1000.0;
scaleFactors[95] = 1000.0;
scaleFactors[94] = 1000.0;
scaleFactors[93] = 1000.0;
scaleFactors[92] = 1000.0;
scaleFactors[91] = 1000.0;
scaleFactors[90] = 1000.0;
scaleFactors[89] = 1000.0;
scaleFactors[88] = 1000.0;
scaleFactors[87] = 1000.0;
scaleFactors[86] = 1000.0;
scaleFactors[85] = 1000.0;
scaleFactors[84] = 1000.0;
scaleFactors[83] = 1000.0;
scaleFactors[82] = 1000.0;
scaleFactors[81] = 1000.0;
scaleFactors[80] = 1000.0;
scaleFactors[79] = 1000.0;
scaleFactors[78] = 1000.0;
scaleFactors[77] = 1000.0;
scaleFactors[76] = 1000.0;
scaleFactors[75] = 1000.0;
scaleFactors[74] = 1000.0;
scaleFactors[73] = 1000.0;
scaleFactors[72] = 1000.0;
scaleFactors[71] = 1000.0;
scaleFactors[70] = 1000.0;
scaleFactors[69] = 1000.0;
scaleFactors[68] = 1000.0;
scaleFactors[67] = 1000.0;
scaleFactors[66] = 1000.0;
scaleFactors[65] = 1000.0;
scaleFactors[64] = 1000.0;
scaleFactors[63] = 1000.0;
scaleFactors[62] = 1000.0;
scaleFactors[61] = 1000.0;
scaleFactors[60] = 1000.0;
scaleFactors[59] = 1000.0;
scaleFactors[58] = 1000.0;
scaleFactors[57] = 1000.0;
scaleFactors[56] = 1000.0;
scaleFactors[55] = 1000.0;
scaleFactors[54] = 1000.0;
scaleFactors[53] = 1000.0;
scaleFactors[52] = 1000.0;
scaleFactors[51] = 1000.0;
scaleFactors[50] = 1000.0;
scaleFactors[49] = 1000.0;
scaleFactors[48] = 1000.0;
scaleFactors[47] = 1000.0;
scaleFactors[46] = 1000.0;
scaleFactors[45] = 1000.0;
scaleFactors[44] = 1000.0;
scaleFactors[43] = 1000.0;
scaleFactors[42] = 1000.0;
scaleFactors[41] = 1000.0;
scaleFactors[40] = 1000.0;
scaleFactors[39] = 1000.0;
scaleFactors[38] = 1000.0;
scaleFactors[37] = 1000.0;
scaleFactors[36] = 1000.0;
scaleFactors[35] = 1000.0;
scaleFactors[34] = 1000.0;
scaleFactors[33] = 1000.0;
scaleFactors[32] = 1000.0;
scaleFactors[31] = 1000.0;
scaleFactors[30] = 1000.0;
scaleFactors[29] = 1000.0;
scaleFactors[28] = 1000.0;
scaleFactors[27] = 1000.0;
scaleFactors[26] = 1000.0;
scaleFactors[25] = 1000.0;
scaleFactors[24] = 1000.0;
scaleFactors[23] = 1000.0;
scaleFactors[22] = 1000.0;
scaleFactors[21] = 1000.0;
scaleFactors[20] = 1000.0;
scaleFactors[19] = 1000.0;
scaleFactors[18] = 1000.0;
scaleFactors[17] = 1000.0;
scaleFactors[16] = 1000.0;
scaleFactors[15] = 1000.0;
scaleFactors[14] = 1000.0;
scaleFactors[13] = 1000.0;
scaleFactors[12] = 1000.0;
scaleFactors[11] = 1000.0;
scaleFactors[10] = 1000.0;
scaleFactors[9] = 1000.0;
scaleFactors[8] = 1000.0;
scaleFactors[7] = 1000.0;
scaleFactors[6] = 1000.0;
scaleFactors[5] = 1000.0;
scaleFactors[4] = 1000.0;
scaleFactors[3] = 1000.0;
scaleFactors[2] = 1000.0;
scaleFactors[1] = 1000.0;
scaleFactors[0] = 1000.0;

return scaleFactors[scale];
endfunction