../../../../parameters/WiFi/Macros.bsv