// generated by compute-ber.py
// table for rate 4 (exact)
// (computed without odd hints)

import Real::*;

function data_t get_ber_r4_log(Bit#(8) hint)
      provisos (RealLiteral#(data_t), Arith#(data_t));
   case (hint) matches
       0: return -1.000000000000000;
       1: return -1.298056274923845;
       2: return -1.706577402482961;
       3: return -2.032113619116682;
       4: return -2.622337485799181;
       5: return -2.955349282566963;
       6: return -3.696359100762435;
       7: return -3.998115929320580;
       8: return -4.874495375914921;
       9: return -5.118258331296635;
      10: return -6.114813220955313;
      11: return -6.320240447391237;
      12: return -7.404732676702003;
      13: return -7.445761333963383;
      14: return -8.699371729985121;
      15: return -8.584570876303410;
      16: return -10.055469071291109;
      17: return -9.778520430198967;
      18: return -11.394016054285931;
      19: return -10.996813409862888;
      20: return -12.742033838208309;
      21: return -12.318164076742942;
      22: return -14.106357550897345;
      23: return -13.366462010909585;
      24: return -15.478777940377544;
      25: return -14.904257605843602;
      26: return -16.976929222256828;
      27: return -15.394851928000625;
      28: return -18.342921260177430;
      29: return -17.395036181850660;
      30: return -19.788979708376690;
      31: return -18.334163665064189;
      32: return -21.365951013303494;
      33: return -19.243738820570250;
      34: return -21.782586334399483;
      35: return -63.000000000000000;
      36: return -24.974956238251000;
      37: return -63.000000000000000;
      38: return -25.502062448741427;
      39: return -63.000000000000000;
      40: return -26.608207634719630;
      41: return -63.000000000000000;
      42: return -63.000000000000000;
      43: return -63.000000000000000;
      44: return -63.000000000000000;
      45: return -63.000000000000000;
      46: return -63.000000000000000;
      47: return -63.000000000000000;
      48: return -63.000000000000000;
      49: return -63.000000000000000;
      50: return -63.000000000000000;
      51: return -63.000000000000000;
      52: return -63.000000000000000;
      53: return -63.000000000000000;
      54: return -63.000000000000000;
      55: return -63.000000000000000;
      56: return -63.000000000000000;
      57: return -63.000000000000000;
      58: return -63.000000000000000;
      59: return -63.000000000000000;
      60: return -63.000000000000000;
      61: return -63.000000000000000;
      62: return -63.000000000000000;
      63: return -63.000000000000000;
      default: return -63;
   endcase
endfunction
