import ComplexLibrary::*;
import CORDIC::*;
import EHRReg::*;
import FixedPointLibrary::*;
import FPComplex::*;
import LibraryFunctions::*;
import RandomGen::*;
import VectorLibrary::*;
import Pipelines::*;
import Pipeline2::*;
export ComplexLibrary::*;
export CORDIC::*;
export EHRReg::*;
export FixedPointLibrary::*;
export FPComplex::*;
export LibraryFunctions::*;
export RandomGen::*;
export VectorLibrary::*;
export Pipelines::*;
export Pipeline2::*;
