// total ber: 0.004892
// a = 0.364000 b = 0.000000
// generated by compute-ber.py
// table for rate 5 (curve fit)
// (computed without odd hints)
import Real::*;

function data_t get_ber_r0_log(Bit#(8) hint)
      provisos (RealLiteral#(data_t), Arith#(data_t));
   case (hint) matches
       0: return 0.500000000000000;
       1: return 0.409991624771120;
       2: return 0.325633766997562;
       3: return 0.251241852472304;
       4: return 0.189079877287189;
       5: return 0.139433872961650;
       6: return 0.101196523931332;
       7: return 0.072560962093229;
       8: return 0.051563538217837;
       9: return 0.036403770617844;
      10: return 0.025580788312008;
      11: return 0.017915695187633;
      12: return 0.012517884549183;
      13: return 0.008731917710034;
      14: return 0.006083941475421;
      15: return 0.004235539640843;
      16: return 0.002947047672409;
      17: return 0.002049720525648;
      18: return 0.001425224062670;
      19: return 0.000990806502318;
      20: return 0.000688710914073;
      21: return 0.000478679735730;
      22: return 0.000332678921018;
      23: return 0.000231199120359;
      24: return 0.000160669566743;
      25: return 0.000111653340630;
      26: return 0.000077589566466;
      27: return 0.000053917582946;
      28: return 0.000037467469998;
      29: return 0.000026036112627;
      30: return 0.000018092409133;
      31: return 0.000012572325199;
      32: return 0.000008736431591;
      33: return 0.000006070885568;
      34: return 0.000004218612740;
      35: return 0.000002931480620;
      36: return 0.000002037061892;
      37: return 0.000001415537252;
      38: return 0.000000983644797;
      39: return 0.000000683526313;
      40: return 0.000000474976516;
      41: return 0.000000330057046;
      42: return 0.000000229353758;
      43: return 0.000000159375918;
      44: return 0.000000110748928;
      45: return 0.000000076958457;
      46: return 0.000000053477756;
      47: return 0.000000037161222;
      48: return 0.000000025823006;
      49: return 0.000000017944180;
      50: return 0.000000012469253;
      51: return 0.000000008664774;
      52: return 0.000000006021075;
      53: return 0.000000004183992;
      54: return 0.000000002907419;
      55: return 0.000000002020340;
      56: return 0.000000001403917;
      57: return 0.000000000975569;
      58: return 0.000000000677914;
      59: return 0.000000000471077;
      60: return 0.000000000327347;
      61: return 0.000000000227471;
      62: return 0.000000000158067;
      63: return 0.000000000109840;
      default: return 0;
  endcase
endfunction
