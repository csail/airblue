// generated by compute-ber.py
// table for rate 0
// (computed without odd hints)

function BitErrorRate getBER_R0(SoftPhyHints hint);
   case (hint) matches
       0: return -1.4860717005;
       1: return -1.8898667475;
       2: return -2.3406256703;
       3: return -2.8292731124;
       4: return -3.3469213830;
       5: return -3.8858839175;
       6: return -4.4400470142;
       7: return -5.0048189368;
       8: return -5.5768836763;
       9: return -6.1539095864;
      10: return -6.7342865191;
      11: return -7.3169160097;
      12: return -7.9010547632;
      13: return -8.4862025571;
      14: return -9.0720239787;
      15: return -9.6582946720;
      16: return -10.2448648098;
      17: return -10.8316344444;
      18: return -11.4185369501;
      19: return -12.0055279350;
      20: return -12.5925778311;
      21: return -13.1796669478;
      22: return -13.7667821748;
      23: return -14.3539147832;
      24: return -14.9410589623;
      25: return -15.5282108435;
      26: return -16.1153678517;
      27: return -16.7025282728;
      28: return -17.2896909658;
      29: return -17.8768551709;
      30: return -18.4640203827;
      31: return -19.0511862645;
      32: return -19.6383525924;
      33: return -20.2255192171;
      34: return -20.8126860395;
      35: return -21.3998529934;
      36: return -21.9870200349;
      37: return -22.5741871347;
      38: return -23.1613542732;
      39: return -23.7485214376;
      40: return -24.3356886192;
      41: return -24.9228558123;
      42: return -25.5100230129;
      43: return -26.0971902186;
      44: return -26.6843574277;
      45: return -27.2715246391;
      46: return -27.8586918519;
      47: return -28.4458590658;
      48: return -29.0330262803;
      49: return -29.6201934952;
      50: return -30.2073607104;
      51: return -30.7945279259;
      52: return -31.3816951414;
      53: return -31.9688623571;
      default: return -63;
   endcase
endfunction
